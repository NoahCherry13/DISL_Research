`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
yJwZLtirp1Kx12tbU1x3K8Diza3/B4lxqHzBwJxI49AqVEgM84pqC5eldHRIIt683xP5LS5+ha1E
xa+mn+TGU3pRAM/+CCpQw+LIiwkwxqhAPj254SxRWDJ9+48LHUFHsdRDPI7U63t44C38H2Oakr/3
Td3lMwE+4iadptaWP6gPQjUFG/8angd0yLEP1lfyuu+Jomn05/5sf0F7GZnBLONRP6iQ1sNl127X
hB49/Y7p9fsYjlcKfTfoGAY7menD2oWLawQivO3SkixDrQ0o8mpAniN2mk4aHlTrtSJ6pjHNa4PJ
YOxyMY6jvjxaRrjwfqYRhWGVuFdD9qTFWVL1aQ==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
AD3MFEpcu2jPEfflXzUk0wAHgOewRC087UMVoTrCCQB2+Lx6RFzgcN9mw2dis3nLszkDemdUN3eT
ztiROlbLk18AcE+8TS54f7auKRoJwkFFsTrs2LfH/qOGFtUn/rozD7nEb28IZ3R5ZHeIiwzL/BRY
cRw1dHUKXWWLHdVa9U1eIvCC99/FPYJqqk5nLTTgaracuq6RPS3vlyEe39GOUz7AWrE2HUphkkWn
/dA41yF+RRkPbpaQ7IfNeQOLQFIUxT6hj2VKYwx1c7xtkjtCV7FDE1HTsz4V3qGodl2jNxQpK+J7
d/9Ku1zBSRFC0OAmY+NlOMmtjdFX+FBxxnFyLAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
iOEM/UK1ppJBTW11F81e9zC0AlWu67EdelR5ygXnIxI8vApQgcY25bYp18BzhP2CpIAiHNcjNoh2
D/e3Mg2v8g==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Aisyk11a+UAKaFI89C72k8PyHf7V445ALAPvYBZylwt+ZNnsUqxOewWZ6z10+PUtmClNrr8IL9VL
CdSiKyx3VIBmXFYEjkedKiWrqi/SwFYP1Nwy2l5FKXu5CsyvkQxpTkeFy/5f9foU8tMueTFrt5kz
Sx7WXIhC0/IKjoVMdIhFode6JDdka8eN5CxXSsIVAV2ekiTjhUQjQgGsed7f8tfl+SXCEeL0cE7Z
GokQkG9H31Vre0MgolLopGz1KrKAo6E13TviNHvKRyJ3RR86m/6XjBw3MHVu5r5NtOmD7LJMKqkJ
uNJFuEp/GWxbni2AkzAEv+jYwtDPe+vL0YJT4A==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ixNAzYel4pLqUX2CEuTZRPyLzeWwzFYV7QAlC1140EjeWFZQVpbEQmFJsXOvqUsaSXt7jRyKdkVg
kDd5JYIogH4vBbx0CN9zgV+RBSNZ/YUfnfeXx85HIIoqmSC/seVOaerN0MQ9yH6PzckoY43RQBXR
xmm4sgt3IWA6iBwyVew+9ACVRYuTNhvhpV+qo3rrAwdtOJo/DUCmsFBZt4ThaAzG+8V55vj+fW71
hbleh4B+WWKc7/A4SJFOFdjc+MJuHIJTFf0mHIfoDa7H758T7+TYemDkerKujHAekqP9MnVMun+p
TF+DYBGCzL3i24QYDah+9Avh0Fm8YAi/vAv4mA==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
SdS+XbKiu+3DB+FGlXKE2sQ4HIHOS8XuEtSHSklRho6GhTYcUgjIE+2QwL9GywqinJrrtZxhydTx
8JdHCUtaIXYRPFbI8lCB1w5S2h+MszXy92ZumUG7aU/ujUIXHoflJOltdIPL1ZA1x84SaMJFMmNT
6o5W3lsbHTGyflvG7wQ=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
pI8dOzpmcrX7Kqik0p2S+qPUFt1/mh0jOMuhSCaWImMiihqw2Oufk52sq2Z86wqQ46KKCipETEcD
TGYUe+h7+y0gZUawxAdxDM5ig/6PcY9jsBXg99x8cKIertvAfzatL34ek3NGr2+w1KrCwQ9w6rvj
/wYTQ4EXd0U1wYCJ7j2dJ4NF5vkA9jLJZdsWVCx9laeJx1DBPqH/rS0MJfThy60PVOBalrTLFF8p
t73RE5lIRnfWvGsDLGs0uGzP8fEF8GVQk6IayAs7Dwmh+thbHRTO6t3UfWYepufFxRc+Sa4a86xz
Gas5f/zDRSn5fdDlricx0TmVLoHuMiEMuHe6Ig==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
MuHeHiXbC09coAz+8UZ1n5Wr1HedzgTG+wykOa/jhpbr6EzVytOfTMGrldZiz9jDyEdgc3Y7FyLa
t7HvsAdHm9WRSIkCbk0YR+JIWs+p6fFQUh1Lz1KAy/+ShCAUYgIQje3paXhCnH8KsY8c8HqHO3YU
DlLXW1n2OXXchynCh33vZdn22BTbQ8lq/O5qbyxcN9ymEkHYjfRGE3C1ywWZlzuCSqNGzt88Pzll
zdAkS3Mn7V/ewCr+ISi6FtPd3T/KAe/YiL9rJV5p3/VhVDc4Ace9NKVO5dlljm64J0h9zE3yWOwT
8TLaEZ6aK1uNRb1IbQV8LbHvlcSQdwxd9yJLmQ==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
BDa2L45Ujd6g8ZEgEyuposGK2RhCiJQpOuKzsQCnLTSBkTlgXrp2e2JnDbVMYS8p+ydZOpPlZsqy
8CDG6obPvMhbtxu/isCJHujoXasvmYLJLlrHRAJgdSxSHWP/vzztRYneVaoW5FPeoO3q2t+45t2Y
iV02T6l6Q/0AjWwnvaI=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_01", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
D2eArKeuKsHAGjV4XokdCvMjukRziARWLskv7UpLg64RYGFewsWhCo9s7g0jA6472zkSrlV/vLUz
WdXZgJjIab+GuMmzz9nwmUrThWiE+A0RLhJrGgJcovtufGRBvVjcnoZSExsERg/wZWbFTszVBu2J
bYnIoYGZx/ypKQIBnRkSVOnIJE6NjSRAiNtv1uYK6cIVi09zAv8R4qxW6vJVeG2tEFSLVwJ912cw
mXmn9+lvHZTY/S9b9GG9bU8Bvsx9GhO9otyMW48aOArQOiM+KDVpQHprES+gTDbMIXcjR2rVXGkR
fxoyDdKN3OUe2a+oAAFSbWwWmJW8VkJ2sx3l+w==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20640)
`pragma protect data_block
NfeyxhwOogyoa9r7frjuqkE4xL69TVf3RmPu+iLU9SF6KoF0a/H9u4kIeOEHNcOONbQFzvrPs45r
dY7tQoUEVgkvjLCG84AXBTL5EdD5yE/u6Nz19Ot0mA1RPKIBfW+zAdPwEuVmF3OJKrLAisNhbV6B
aQ6g2AWMogEeMkZUPC2oiFu1hTsLi6VxMHtRvPS28nmASna+KY3vgOuGSxIFhn6GFhP1q1JYn0Z1
HpjhmqepU+F0jmDRivF+bVY1k55LosZJ64YjSM6VMMlDVvPaBdyxbdMhsd4mb+RjqNuc0KeYMG26
nxhg1JdC1Xj6kR/ewGawF5aoCAo+w0nzslaMxxgdFeYV/aZMGoI9V2i4Qy5JQwfrUxPTlCON0jrV
Lw31dqzq8re7OA8EfY4elmAnwUThiH6iaK+TjGQUW9irwzxFvE8/rmjGu9F434x9URh5IylZ1Kal
vhH0REj7IQOtXhjNe4AWBNw+DkPgnOTTLAuSo0jnyvZcAQa5EBS4N2xcjDcpQbHj9cPoB1tPbY/Z
Bjq3iERsuZrHNGtDKD+SOOZHa3j+R0tb5pj0r1p95C7hc74W9ltz8SsCKHTRH5Pb9piQGafPHbwV
ywF5o40RbmHLl1wISdjNCKH2lBccuT3Q7xL8pwKLOVkGDUWE7Z/WV3DE7hRI4J8KMPZKOxEIxYeN
zYEIrvgTwkcXeumjK+CcdapzAX4CgYSxTXtS5p/sDkhHzlE8CS33SR09517MmXfGVMK2MYf9AUWR
iBlGMppUuNewCXdX02aDgIeGOhncEzdDgIbHB0V+QwxDTGhw/PLMDZa+SSziqmmcIJnPYLa3QC+L
SMrx+0C4pVG0cPhHiMHAQKQebC1SAZyUwRHKM9TQbeNwGA2REyuOYDE1PWOfNSd7AY3mZpHXNiRE
fgrAMXs05ANA4J6ZUkDAwHjpV3lU9ArZHYw5UUm3GrqQXbG67NjKclO2xfTlvMRyff5PiiwgVcXr
hG+ijNixgaGV+h4mjUy48UESdlcpMyW/8xyKo/03qu8bWZBo83A2AVMKxq1Vw4p1QSY0eejF2sc1
kiSIoUhnP8X2AtPZ7oJeC/kJE9r8RTvUBk1241NrZG24fxe+zP5CKRzSiV9EA00voPu6DRoFu9er
/1WYmngnZBBuBFQju/2knPfIX5GJbJ6yqsPlm9wlIYNfmRFHr0omvIIyVuuW8f9wHf3I8xGQq4CX
F9/hcTQa0qPqt8S/SjKOeYBW27FjTS0ALgICbCh5wlv8J5PtLNkEPHLtH1tMbNUXNRTVluSYVfyN
DLYTjMbRDGypegNJij26moPVYs/KZLd4uJMYPBMb1pW5CH8k7tLBy+Nv1yAao/qS7GmEKPkfQ9RD
S1vtCEmoA/TVl+rf87F41wrPuGHHbWkLpKCEASph5wjsixmVIhAQ/NXlFyByR/AuScujxI/fUmkn
bYFd6DJClWEWxoVYNa9WI6dzn7ZcFf/bjR5fUXIMCwSd6EZGBAqnqwkhnZIqksszdFuyQ2WBGFBw
u23vLoBWIz5h667+sDVHSyjjDJmS0jOOiawDoNNTNd0s84GWOcTidGR+55LNB/goIJHIEO4IEvx3
E7OHu0i71eJ/n1tlnefM1GGKdfU7RYRi8NmdEEtbmN2j6bZka18sLCgD6ylKtPqS6lFK5heccnSE
yc3IndpWT+zy0eBlvC4svqD/Fs4fjMpCwd70+I040q5TqaB/8KbpqhQhunVkyLfQSN6TuNx/vQkA
cdRt6RTxC+QCbfnJIk5kOYTGQ9bVZm3PtUzE5f/eyZ3ocT+Lf2b6D+cDYEeegFGkJbSY2hWw2Bwy
6TpzT/s1eF543H/xB9li/9I9+RDLJfBpXs+FanlxIN4c69xv0u+pipx7iWyN1XiDRQ4mL0dZRl6H
zDfOKlTycxkfsGuunrjmcORfFuoaToWgyDHy5nf4JHKksG6Oz4bFvMngssQ9b/cUXE4LEswxH1aS
Dg0xC1HeFmvhlvlsKSiVE5Z0UxVi4aVJcr16K3MyoGdHqLuPXaeWFAYMRvTyQIgdG09rSMdSfz4m
kdxVpKWGTiGF4SFjlsnoyO6bNXpY/f1rcY/8+adq6zx6y3n7/v8ypkIEsAWuU4WWm3MEngiNJMNa
/Vf4uoau486Em0i4Xj6W39ch32ixtw1iCVukvx5HiV2qMbg7W2QMbvB08Yu5WS5zaHAskCACIIrv
I4SoLWUEnvXwtk4w4VO3L7LwjJvJEofdN7rxh42Hl/IOBWMK8OKbkkza1cAqyVyRIzb1Jvs6ttY4
zVAYi6Ji6lbgEFmYhPqGXCjE7r3FxGsa4scGDl5BNLWqaFAYS7BIgp+ZjstWVVGFsUJs7rkKUTST
BzsPF8GpXEeEPfmfSiTP7bNydZe0SOlxkOibDWVq2bAopyMASNiUwPOVUdqduChoEnRRD26El3gm
sag6lUC+y+nL2Iq0trNka1eHspWrJh0u0SS/aJ2N/1QDgAoh50vf8p64mCFPZUQNlvRivpVCN7iF
tf9lGcdTh+1dRS9T5wxRInn3r1ZuM8s3QBS6BZTTgXa47GhBPN+9+ntMj5Gp4CwPP4uZaldPT4dM
u56dtX8bEUYPn3JW6o1M7cJdfGrJLskU+y8G4NQzcKipeypkCD1BrMs8j+nVEm0fwJEA5AjUUJW3
CnheRO41vIDheB0H2LGX80fvFO5YW1EGTxeekJ2UF90jyEXAKdWjj/ZZdND2WH4/oIp9RQKv3MsC
qowuvYny/VCyyym5Krjq8dVosPDWh3r2Mppq+NNj6Md42XXTqZNL2hibsXpKM34qGizMWJ8tfp9g
BxgIkrMFeaLUTuYc8+u5aDWQAP92GtJpsZmEVLLwqjSNGk7MTC/7gTIm3Z5w9fv6xqvmI70WtN+J
XJ00nicCfyzV+i8wCAdGBldCCkKnirIUunlneEwz164YVg9/lbkl4LvN4oTcUo/UeIwcmnPieH+z
XwCokdMO51UMdL6YqPkDK3TFXKSDKWzANlFJAxUtCouYObMYB0z5FaWuaWIMlREehTuC86n3i/wQ
WItSxfPB38Ti7i8CpKIC/av+oiEGToYb/hroVgnk4VOclQGwWoKu+nIUMpjLD+E2YpyKhw5M5hTN
0nWx9j9FkQ97lPtbfCN0G1sUbQpoY0/ZSxK2Mh63eHA1abHH18N76WD6CK4wMIYJIH0N+sLbATEC
GCD8PcZAHfBEt1spmelydgO2QpDOSNOeIrBwLcD8eCy5t7PC+lynRWM7Dp8InyjF7CoozPz7Zsrt
UeD/PkFYKm0dP9njnXkzZ/kWATQYU3jWcPMl0UCr/PKIsKma1C8VHVGnIoFqssOZt9H3+XFMaMwy
cmNVgacjYWmUk2ibYsjJULHPUu4QS2TNswoFASEoEyHsoqLG3XTwIkHdr6L4hq7XLNSUh1dpgYBx
iNgEqe92bQ4y+DWQB6aarypj4fKDFKJ7F0RI6L4PJJQrt+EEYMDwuS4p2A+ZzSEjbAjgrqMYJZ9W
/ZtJ3bVeiqc92lL08/Q7duyeLi27LYBwKoAEuq50UAC+Ad28YLUJuyqZJdw36VDrsP34RAmTlJee
fDarbDco6izv63Oon6SzAtsRXefyRm3/SXOsNB9Mb6ww3C1gCdpVOsJz03WFrHKrTmFlf4QsC+vI
4y2VhW7nQ9tqAWBs3BLyd35Xew2SfrKTjf0B5jAWvGEhY2av2PcDwlvcN1TwpnNt2Ino18+aSm4+
Ng43XU67p4ld4bEl+Ek1Xx6bBoNNIV/dbI5XeYW3oWHaV1Ua5xXPMfsJo96KIdD/z81fqlOoI153
OFkkPoOq0r/TIxrAX00bhNJ7K+khdgKJRTKYljy8oJWXjkdx8ApIsd/L3Whh94G6qdcwwRvWHY+w
lZRSZE0s3gIDXl4c7NMF3NxVJHTn3EygKuifxbVopMe/rl2oJgNjiJQ3fQk+tXbAujVAi5bpOvPW
jGk7/oXIRIGLlRVLAl0jjXe4zinAquMLg03+a/59ND5Hua1t+9C/pqqmwC86rcHzF/cBOK4vYZJK
EgjNVk4+8Ni78+LNKiJYe6mu1qR35rGcJ2EJYQ2X8C1QO7rcBnzIXO2fNGFZNbHmlczaBFjwD4xb
AFIPsAceJAYqxqpTpDiSVi8dYqwLpTNQn0WYmnZ1kS1a7ZfGezbFa1Y+KfiF0c63xbNzxc7Dox54
q86zdV4x8JlecrTY3V33AT5o8rKy7Mr2D19HB4T0k7/pcG9dfdwBUa0t4k3F4V5p953ZZpkCvNlh
aniuf17018Z+xHbs51APp2YYjH8StgW69+iVEKLQ/nHvydmBu+f1hkCcZHhfoEDVj1ahQBbJocjW
c53WN4+Ch15iwL6x5cFU0OGERnjEYt/cPlh+TQzpcSxzA9+YKqkYJnC35vTjM3A6f6hZhDlImbnn
ZzANWHhncjKGamQRW0hfpjBSD6GLNgoRKnttfuPhbiAvrO2pr/YlM0gxh9J6SAzKc8JxmwcR2T0m
RV2JIrOHn4BR9CvlWD7nZ+lS7VoSIU7q4dj0tdVM8gzn2zIyMw87DXg1s80OMKkfnEKdHK72b6xM
RUfGWLZd5NVq03efYdx0zAe/ueEzKSEBCXaR+1d/f8ftDvriDnqm/xcW3FgqZlLMJke+7JOX/KBW
Z7SR1yhqDJus0DhiPEBD1rXiWzYqoaijpsLXsZzPEQ53A0m9FpofuoLUUBldHHX/ZD8pPaCm57N1
S81wi5aF5cyK0r5hKccg2nLVBd/S4YnGXJfqP+RsPwQ4gdsrbYDICBS+1abGfLU4+fzMEcHEUhv8
S+BpAMW97mQnjuKxu+Tth9TcxCou4rOeNbKNx8Zkbi5b6SCafGbdhTlSsHS4hwh/Qvd+LzfD4hAU
kjHVDH1r/w9L4nl18mrnXrz044GsPK2AlF7prrlH5BIgoAPIovtkTCnfwRFlNYfuOzSOwnCmzWyK
tij6QVK9+O2rARYIB17kWBzw3i/7VYfE9jNfpqFjazzoQP2dQuL4cbckZ/eOycDPfyQKnOLhncMO
xvQ1wlzZoOM+qR6LSPrt1OUGoLTbXyZNCn55aMbVBDv4dHdZCh/pxDs6uGOOal7NPbJLy8x643VV
gHKWj2JqzRZTih1W/1BY2c6NHIkG6BW/g7VKdnCfP4MHyN1RwUBKav1mOgy3mEbSqg13IgOOs4FL
qGZdkcw6aD7/lvv1i6m6qeym9KvbsGFRTkQ81X+w57Lhoq+zO1RYhTe97JiXut4ruMj5qTU3CzKi
b9Ci+v1gXLNE/M+3vtJ/uJsdy2nKyhfSbormJsJ+SGkyGCQslQ/Gy9vPc/hRVjQIJqwC/WSuKud6
fk81m1ZgtvGmkK1NNukTJhi5Yug8p9zmQCSihkpRyIZ3b+lJ7FVLup6pwbIHwsXUXQBY/dSY3jWS
gnZ6zXtkhB92gO3bYaYwvh+hkh70zD0t9QkV2Un8BMg9M+QF0J3pr9FjJCSp9afp58Bm6YA362Z7
N4COpef5qOsygCF7wixnoNXkkpZgKpi/QGfankj5yXrcaN7eosb1jDsTkPd82oR4QEqaZZ98Y1UF
1vKRC0oDvpPwkqtC59bLTYfdeB8X+FiyhtPV159aGyYBz54FIYtcJARRekTtijuBiCX23Gt+25ZD
koeBSpD3RCY7kWYujY3RiMcZIo7Bz9Kwjf4bF7S1zPm010/Np61c+ivUrsqH/+xf9KFc4PBWGZMw
pm3p9EWpD/dIdFrAWnkKok/djYA4TMITlIBxAtttdmt3OJQDio8aZvMWpRwBBK4TdV4ieA2vq8OR
CZts/HXJYJEwJYP3sXfspedpnQ2LzK9/rwhDvJLMWyfY1dTYV6b2DkKCu5BsXhXjKWTH020HR9hu
bMVpXVgi0y1ZMnbrsUe4WVUHDx6RbyG0fL3/IKkOZVXTDPDS7cAg4v53+ipO+5you8sRLPiCaLfS
ZpvJSp7Cp6Ta6HVMfI2JtBtZPOk1Wiibw9cHBF10vAQsYp107CACsaxtQcnvANgD49JuK3pc7vYq
v+/sYlgd3Fx96Oc2BwlCMpTydg9mDfZhxcNJUNNVeCSjVnLPTW2n0hMUwoYl7lxXxXY5nkeQPjwf
9G99hXYNfepPTgyUy5333ndSMhwc/chvTLEbWfCqqheWc5pg74sKFXhLRnyaTWqzzgR4iA8w7dPA
kj4enLx4SSHD6sOkh9f0HyPrHg4tHHHys3QLW6WxFss6f2Re2wdRrXUCE1wAfF7V7KobvxBGD99F
ZyW/45x1g3BgbKhOCm3qTqfSkhM249Yzk/YQ4Yk3XXX0X632X71euDPKlQ7KhlDDxu5XFNoanqi6
JnO/GuwszYwROc5VzVD+1NrQaMzmSrV2c0ATXDGU2SuJiD8Vl0EnFlIi3/3VsSUPGmH16eaRBTUS
kphvaJrW84wffFyL6dp9Jpf5IVdvf7xahzOyXWMzhGK+hS16nKUNEYI87sZ0KCLflg9BD/GJSZLm
5DExAUhy1Rv1fMdwLAApAeqlH6lD6Gmyl/jlsYTNr+8FdvXTKMWTsRZ0KNYUWd4HKns6BZqjITuy
Y5h1ONeJVopxbLEhr14mx1g4hGKWgJPG4uShHwDsjRmOddz6PAoFfAdkthCSNaAxm/c7zbeM8Mdl
5QECQC6m9Ko5PibwVWlDPWs3jq5QQZTwg86cXXDHvTpSNdCewLhdrKfOzv9kREkfJ6ntkS86vbxv
PJIHYcnSKUXUsGiWJfHTFACAvwFFImd2mBSNUAnPQ0xrzISk1TFt/KnxjAX0pgTFegZ134W36oJ9
Mli1vrhBmCvPn/P5aWgPWaBpIClAXnQtSDzzyxLAhXn6WmknmxbbFiTJRpp/gSKOJkCwihuNW4t7
NTP+V6+O6F8fhi8qnMlP/CdbRzRPR3Cm8b6KxgRPSY7IBbs4/m8Wwzo0gkHf7AhNiA65V96+4PYY
eVMrizF3aICYGkhsrVmBNClWR+fkvKb/pICH3HvQCqIXDrVwqmKrZh3qaU8Orh6+bQgXEFeqav1R
4rQl5EqOP32cqIkJV/NuQkgkf1RFpiNX7YXfhuBJI15uohvlTd+kbN8abXQTVz9fV3YZDhZDpM8M
qz6CPIHHIedKmTK3Kd8kGM8ZDkejfyC5evNkTwVBJG7Rd70NPCeFS8mX0X6YpzsezEApzFF6pLvR
4uObFHGmjIjPbbLuc9YFysUb0IYBrfEwdFeXwRJuwYU++jw+nggd7GWJCjd76IgZhtUkqxc7nU5Z
oCYs6HB5GYVbtItzFislnbtWzu/7JZ9JB1nSujays2gXVx3FyGPateRYeNm2V9eNzeFFqIdO+9Yo
OTx+VzGqD7pacQy9oe9iGGuy8Yi60BPkqO0+0dhkjg2ddoPY6v3rV0FzFzwlSdORORsCveain6fJ
c3DcAgXfVnxPOGPRtOdm88Muro2wHzQVOOJxNaJwbJ/urwYEhilupBZDOX3xcwr03v1SJpnWEcPQ
0Jy1cIuq2Dnl0QbjYMOMFex5BCkWhtXrraox6NCjkClXHqnRgH2TluqUw6WLTGdakpG01a1I2kUK
ni87fFN4/r1VT0EP7XZazf0iOeZLLBxeiY3TYlZ9YerNM3Iwd4OjDstB+ybjfrAbY3UrJuXztYG2
Y4+jNg+BknOscf3EpzJgboWI0YYYK8Wo9iDgRHmTkyTaAqOi1EwHzSF40mhvwFloLYZoLQF55MkD
IP6E1J+8qMALCaWUFf10sYNvJrzZYN0/fvW2ewXY3/0B/axT7lRF/lWWriYlEm2IGC2/RjUB0r2f
YrpeWsvhSiXcoLxQ28U6fpqK+Df0PLGOE16Yr5/yao2rMjn5ggXdSh8jji9JpQPsvwUOQl/6XxS9
Kzl/bgZLbOuAV5wnjwWL5T+zj1WDL4SZsKTw0oZ+Lg9t/Ln4PvfTTfiEFEqnnBlCnU1m1YLsYQvw
Msc7U+MMEyIZzorVyQue7roTW/l1Ecib+KaDfhFVwp15dmK2FEMbymMDmDTd9PNimrscGX5KgWkY
zjzDGGkS9xCaNmP9ZPPIh1ydem/jkbylsBhM9ghpzbWiFUlAfsbXEnYXGmpyGBqKp/BioEXpK6hH
Hjf9lP41zy5Cac74NdVMQB7dLrHInKGy5a516YyGHnaeGxUtiAGWBBLj1byYH/PIjGA2mTRuwUxG
aJCP3eu51YOx4ARCAGkMLSo1R3dQvGPCbXqJoW9SD7lsH0htKAd0eFWc8LrUOeiilauGOpHOul1v
87Qyrxf5MAkM1UIWi6tCv9sFL+SiHVgpQH9NXwsqx/u/WopV+IfRTebKmxkub/9cr9ukIXHRaMYZ
ul0DX+BTTH4GIZ/GXasDuoEcxQaSgilN33FyN72M2jd/KOsxvGcq/X+u9+QBqLE7c4K2QBR7kRIz
qe5lPhlpaLgb4Wfz4XQtzm3glvQ7Ej0fgiqb3H5xyTLk1pA3QHk5OUOfV3W5xhIkAA5JPprGd0Yf
KqWReBZLgS2GuE2hotDkH1qVuVXYs2zzbqby4/Zbk/xPDaeHh3O4tSLwGyRZ6EWIK+Qp4vLnGvxG
WiiLlK0YSE/f8TZ7zSit+6ANip3eOM0bhySGQk3ZaomAW8ilVL8iYSYrVZR90ezq4nZh6WPTMyNV
TTJEvJbyMk9oLJqFn48i3baLgxNeaKnchpCp3aJBezpBeQ48+4pa9uuFeCPsc5CMl4LD8vmH6VUh
p2eAaliqv+KdKiGvKyLEOrDRqNFFFxsahoEvb2mXHtTBanla5HCbq8qhxBMOBWiBmgqiYE5PQaa/
i1tihEAe8Vjs7Ps1ftS2qsc4ZYA7eLutbxwdtucDrH7dXoaS9e72idQpM3Lqk8IDaBFpGi3Rweu/
NiMXfcO+bsDqLvFiDj1xPEofQ14AsExAeEvbYXkrkEn4IhBgV5SR9a9e6VJDnJjp0zLd9C9K+daa
nYl2jyHVBM2O8WyPtojuaiOuYNq1v2STMPadprVciDeqLgWwyyAbgYbYztXOLn07pbJ1RfyrFSZR
0xzQ6DccrPudWmqW5vxLLY+sRNEbM1sR/FrNGPrNVGY+VeOGKOHA67gFo+SqSaPvPyj4Tc4Zxn7C
yXHP0TOQKxHCokw6pPBTm7fm+gGunDp7+Or0i6WxJRUIUl2eSt5ns91Koub5mWxvhsB5Xt1Nwsax
ujak12YG06c8+j2YJGLPVVSuc9kdUlYDoJgtuFMvR1E+j+9qYrPqV7ncQx9aj+/l8xyXl0aTs9IG
kACt6eMo6ijP9Q8QKY1QAAIAz8tyQTJHt6JF2x1Z6uklVwZ1rFj/wpfrlEufUj47OO4Vk+o/gwIO
hhpYEFFHwFbZs/+nRlARYw8hYKxymtrisHCvtQos6pnqjyzElNtTu5uzssRow2Smh1fmvRYzcB/X
zQ9Ry900DvjCqBLaRKCZEp7DS2SRSnrDsETWiVlG1hhS0GqYOzbovIWJQxoIY0TcDnKYHpboz/iV
Z/x2drW/GCNkxUokSA2yURVbo9K1BpyZSI7XteMXpZlZgjVrmrWB6VNnKxaIz8kBm95Jnhe9cdIq
P80MYBGHblUHpZEy3d22e+T+vxef+N0IiRnYNvk9BKHEvm+kLKgcYLwYIIyCemMRPj2ousP78G7F
klwZLROApv24iJjNVIwqD8QaGf0rm/ww09T7XVORDJHp9hcFwBx2WQiVl9nBaz1s5oP6G8STqUqJ
/OvK7sEXMv394/KCvmILIhztVGqFtirJiqTXDHIGKjIeX63SViYiGrjc4p5fS+5hhjUQGX8V+de4
1YqQ7xXHnwol6SayMX6zfH0XOAFSQKZVz+aCZNp5MWtfsN4/5hOGU4zuSR1LPRD3rTtTjlajEG5W
rLBZREIqkO0MpfHG6PAZyShic64dF9Q16NQU2wDgAncAgC8Md4SQqmwtgcG36gpeZ0mN2oqI8FsF
jbKqgZs+OZXFH+n862r5aPDVptQU9K+zTAdc0LmFQo8lDEjppwv20UMu3YswfzIwHxG09stPZErO
b3dGXZhn4lCLU4F33WllrXPeDaE+S1ePcmtPfWyIYk4LpavCXvQ9DVRApK/ywT2OW84tvGrTQAqw
5IS+hv144KATShh5D6EW0NA/oFnO4f/3xu/k8yF0ydnSpeqXJHR/NaKYnDa49otDGvQaOl6xdhtb
u3aw13A7sOGNOFYH/UZuPOWjTiAYi4GTmUYAucIOxd1HSLOjzWEyasF+zmPIAORsQL4G2SUr4suV
3V6uwscn/oKNryuYO5F8NGYU3Ax1R85eZmV6pxnwhWhTvGNjLfZg+TKQbT91N1mYruDsbQKNuNWz
DN3TWQKoKF1abKo1EPV+UtB2jooKtHorNePhSl+BwUtz/yqz8g52ezbTsnG39RuIZImzHl8lJsGU
uTgrhpzJC6tivWsckXRI4KY58rzFdffKc7kfkBQrEeW07By9cf47o4fZ4/f2zoedd/vnImIjKWNL
TA/zs/QHvAgjCd9XPJp8Kd8MGIfbwGIV3BjBZaAOC9tF9O18EQqlSMK1j2aURJ8Stog2ZEK3VJTP
j3ss84iM+tCBkzWBYWclxhTu0sy416nLGy5P4SbJQGeiVbwwR8X0wYWxnJ+9gywtZzXUGXQH8Xsr
ZuE86s8H9oY7QdtdgtDQ4lJHyCdk+MtYMNifMVOJRNKRORC9bl724koVsa6mMVHwq55brl47qYmZ
Budl6Pa/8Nr9pND2v8PW5TRwOVcp+olJLUWlULMi4RDNWfohYy5JRi7jkxgvlck3elUOCdavM36C
lmA35Nt9glGY4flvp+rrZWK9PsRVZ4w9vDOgeX2h15mRPivGkGa+qsmAww5obaUnSCWcU7R2Miw0
Y05vJuqpwYMalvZQ206xdvJPOXv0EBjZkRtPI1VQGPSJeilF+ge/Jd0gZjq219Io7+P0V/PEkYvj
d9AGK+ZbA2y2g0n8wWKOtkD1MowOTNVdHTOsxA8Y7t5sgOf+UwRjclZmsLY97wK2E93qx1OE0IHE
2jqeQk0yHxpnI4InrckhyWh0KJWjmNNST61LndFWnPbMJkA8kzXRbvBqEC3FwQ8s9qeCXFJR4sYA
bs0aYep9HNog1R/PYqBQ0Gb/Y6a0nrZT6BGYkcZlw16yqOP0ZqMqgF75HQp/eWW70MwKWupgZy81
r7XUABQEB3UiayTGcdw64JPJoZU/KeebUoOUR3sg1+GETfN1kaJXM1+1e63sTIx3v55nU+NEfkGV
TMbkX4lLUWb1GgpcZ0SMxIy1df6TbxfM3c3a4BjEsboTc3QtX/mBJWkx1bhlNxe8LKNCT40tjmMu
i6FYvN8Niixq1J9FoMRLRdsHqzDgF50lOjEXxwt5cbXw4Veia+PeXPVkf2ZIOYkC3AsjLuisoNAy
yUh//JBtEdWEMVqhAFbQxixC9Sged1yg+MQsC3532lyK7gtluLZ9pmanTz86V+OigE5KCbPSiKIu
ct6ZdWdrc40RuXmgwQccqYzR83ZR+xzkKVuhrsY+Ofx5d1PwXz6RirxLgXhczqjcx3MtJab8uOks
79LKLgoiH+e19QhA59XnH4Pn385+6wa5RICdHpAOz5QAN6uNzT3/fe5MtwkwsvjuLm4XuXd8lFUR
bBC/GtUq6ztC4eu0Wxtpe1F8qIqniWhyGP8/mHqzm8w/5bKdaAUbkYpt+EYr850kg8qBaYjhrudc
uqlJa5vhVawVAC2rT6mQExGLk/6DUDwQZSvo+mI37ujMYglbBxCbZ15hP+DwgaWL5NlfUjHgjSfX
sfZUk3s7F/JW8vmE3RByTNtN2BuGHUcw8wtRJClw01dwgFsjBTh+PftuCKUjD0/V/GA9k6YFRfl4
Ui3XyrnW5cka9kAraBoukayMIrdT4kIDVxn4EXIiCT3EJXOb8ApsHvyOH4z9TqnCU5wpqLv58a5U
pKm1v/vbnzaIqmxNaYAPnh7pD/0b3f/nXSzwsUj0vMBCQU6ogpCD9bcwqlt/9IvmeaJR2MmTtR8w
NnRiASHp1Idy8hq1qQDdb4ExpI8an1VLPeYvG7AGuD5mQCYFg6sROX1lFko1BQKhvDwPIjcmNslR
Ss0Xar/E5vCRp8BOSk07rxYr5BaUyOa6eAvk6QnXqMyzGcyalC/+cFO49/bqnxvMaMXg7c19HacA
SvZHPSgdSqD0hh3H+1nwXCb5TnX7EotMXm5qRI7LL2/wbo6iSZ/8RpACBLTeUwF4m5tsji8z0jy/
DUJEK0n197cAfLez29MF71pgkTTOhnq1xhgDcuwMu9z9rOF7y4oDLR9EnnHeU9WRkhPJFp/YojjK
8MUCW8fEBOpOJcUp0hz0NLrPwewQ7caXc46so8HJbJOcAGxVO9YDg06OzvseFMh+da4FtzN5wB0k
TXCbn+j1pNDyNYXebxksdQoYaT3XJk2Jue8DKy1hI9L/5ROS+ciSM20aZ7O1G7pwdnGMG1+xaFdJ
lkJkbUdXdjydVWg66TEz1vzRfVVpdG05EC3pWmPaWTJ43STPISc9ekhZQSwDNlV+t4y3rmSYN/rz
nDBrGBZbe0r0XdrCbZNX1M3t1hPN7wYX/TZGj9/DuSQg0fhwb1pNmS48NM1l5ikZ3ds4b6igSO/A
eE8azLVEAwJfPHFcVQ45GhQTf/EL7vK+z/yjphF4liQnMUCxvzQKarXQ/H8cskKTDI1Geo2OKEnD
Ty7xWxDVTewxGqK2E3SX+3u7bVO1hot24UJJexxwvGDkSkqFwKL5wzANYqWFrXAQLba8/oSwqW+o
PAQ4EK7py7ezOvBG483Qp3miq2y/kYJWxJa7t2yVgcEHa96EBbPd+MxMQx4VsBtA/K+vruIsDyWw
R3UY54Rn+im6jt5eyP38/xKD5oDD8DHlC+HCTF/7f1M3HwtbSOXG9QqcpTSspupKlcHqZZRvrKtp
JgZccHe8jKO8FTeBNJ0QdDtKPDVaJXQPXg62KFuuqjAjukZ6DstM3cN1lpMmvQdJy7RQt5j/uHGs
WN8Qa+BO3nvYhcJ3T9SsO5GTjHNytXvQw41ld/5eN+ilP5cGg5J7MeCRQmKWjhhmU1nF5aGA3JaD
bJsPCrgUFEYRn0xAy8Ha2PNbJ0/c8l4zbx6pYXurKBeJKob/WOHMeS32br6MzB5+FWEGw6xPbcu+
dJwdGjpWwP+3+tfMYnaJ9Na+/5hdJ/4auRbepr3c9npge6mCAN+zsqH7l3uVUlw8bJyRZSetafJV
E4uLcwKB88mMhkQQeGOzMNn8v9AnCCvUmm0DbkcXmQpAMvfdm890Cl1a9CvxCDzTHKDDXbI4+Pfy
vZK9SULXyS3dW0+R1PjoPwM2eNRUM42DMfJXDFg19LIRkNZEU1P2Ve2JXGB3kZlQs8fGk+RPFsrW
hp0BEsQvPCkRhbCujYKszDOlFUVoeyuEPO3XHuDIj9VfinjrpNNtJRUzpPRKVWgqeL7PmZWdyoQe
JxiejhKF3LPXygGAai9xe1Hcn0YKukgEc/xm5x/o6Eyl5UzNdV2QeM7CeXpNQRJPNVavY4pO/z0B
4Y8FabVoNiEI0qegvb9FOIF4cFMclmZTmaPPlLo/98M5ziKSJ5I5pQQm+2aOyBZLISOC4WDcPcmg
6wMDNeNIoO+vE8ReeO8NxtjOnsIU60OT9B71LEfTNyAYfPDLvbHa0MdrQo8ffS2w8AlPsJR4h3sQ
K1+x2SjYuGFvLbcAZNQpTJgk+q0ZMwh0pN8cEOWHl5hjMKsAxfuVCGMXD381THQk7UZ6e3mMqXb4
0DVk324eVLvDKdXYjw1WdIWVy834HtrMoUcXK/IveCxFEIZgI+d+80kr6RGnoI3WH3Wzi0RVEScD
KqGHn10dUB6Xtrx/eUWi21gPmDH7sv+C9d22CN1uLASAs12SeOHJSOR0WgYqHwPf9NUUJJ/NBTYx
bZZxKLJuzW141YdZ23oywCJCGE+PI3RvWJ7wZSLovzEcuPsxcVrH9RLw28a5Bjnze3upAlRxAjp9
JK9D40MJn8gaOYLwi8pMEQ7/DD6oeD1DmNO4XAQPNU0d472jGn4VJRQj0nna+X0AWlKDretxM2JU
3rlnTRjnsvy9og38nyjZSIjKSCWKORhFR89TfdXSuRpruQIQwglIh+UxbJXVFhrncygiV1JHhqla
kzSzX/QY4+xhqqIcjIiw3gwWsiUk2U6/uujzqsH9f0kbSxAYNLtO7sxm8QmVNYJ3OTL19lA4q5/2
6PFOX0ZO/VTBqTJ0MaB2yKsEtn10FihEkGYfsXsCgb/ELn5BhPji34WnRG98H5Oq4cyUm6y/5/eE
cMrBbkdiCPN31GmAVjVdGBpKdcQJraI5x0/OjexJgH8OR6CeyTR8lPxboSJTNFzbvqyV4wxhP2fD
wv13InSEhopZjNcGKwls+S8QOGli9NaDPZ5ipXW8BJxZK6QFm5bp1PnhCjbhD/Kwu/n6pUGG8BGH
w8fXNeOTTOWzy75xcTzqY54cE8CPH3En/fraB4QnjGcf+b8S6jYtHT1UwZMShpY4afw064ou2s0E
QBGHnZsDu+jrodIJFc1ZgHHaSYEAWP/gmkdcCqD6Qg3GA0R4C9r+Lt2gTZSXE+0kLBD6UTNNB+0W
W9AEb+grarXI92HCZ8X58F4VFY+HN7HeuSJvF0OnQRLGi/eiw3eH+Aiko9g1kXvyW/tt6iu2iBbj
Vpb8bYIp4aeNyuJ+HQVD6hoNWYp4oIw78yjkwcYCq2sj5ak9403uLq4/pq67SMEdEAqJvugJFiHg
10eEq9gDgp25MpoJV52dXVbzpxbladFseluQ+qilsOba942bbvb8yDbcqHpudIJUIAlelzGJBMTO
iCH71e9v8JnhlsyVcIMUPkkUO49IosxBI0olJjNL+99un50iuVK/bdzqIvcrgSykS377xk44xXSK
otonTrXOtmUXJUaRtFttbA/otqyCgE0kXp7BVz1rPQaD1lw/Fvvu8edhFQmIIntVXqRCqlzv8lX5
4q77W5eBExCJkNEykCpRbgkN9sTNJck16bF4UIonQJlXCCBIpkYFla8aXYzD2wg3URi3QPsY1X3b
wTF4N9H9O1DRSrkU51CtqinEItMfbeAjHsz77PC3PFd1DuYp9Ld0gtdAnXOrENSnYu7AKLcWfEw5
T5r/RQ3EieRTlvBwqkphDZBUS5l6sbTZTQHeze4s9XKdiinbiqYnkqoJWnfUSeDkMg5HPdrYO1df
kQ+6OsrXIkmVuzrEauO4MxIMcLBs/BIBLhjWvZPDe6Pq0yfj/2Co87ASTeRQ4D3Ik1jzjbPO1R6Y
rK1/zNiYCX+RtFAaxMwBO6Kt2HHh9orCCkugwwPvVWefbhI9448VPRQiMpwgKkLt1oAYPhUnUAku
Dvhh26Hg48ENGdG0TIGsRZhSZEZ/zljDFkqLwiKmT55zcllkp5PpDUMDIeEqz4fsqClmtAhZtJ5e
bq26XOWdIH0+EYJfig6VT5qfW9lMXncP54BywwwCW2HNyj6Z/LMYDrISS9QZ0Fh8QQkkNXGGIQcr
omRDcJK9sCg2hPZPufvbXuvqYIma/wgGzZBNKEX4Npy1M0ai2ygdOKJsMCPLSNpwjDwDZwlKHrx4
03PXlOGY6FEF5KZaYDwdwaHBOKfRN64SPvsJCccTbMgi1CGSDeRX2tjcyI4Z8UIDCsGsWeSERGcW
wS3YaqaaypFMuzd6+lLCfOW3aGFL7G6onunWSe5GycvZwlBkO7uVKrJ3u7nvv15RhvhJOFaX9rWU
cDN34PWX63HqVImH+7Z6cMKmxHuhYOZ7cAvN5hzQuvv+n3vkV9v2cR4PuXs3pUiQpyLukkVeZVsq
Nl/+EkIinw2nEieiC8xr7AdTAB/U+QCc0G5daL00i7ATKlJJUiDiEzhbjY5mWArBsKCg6+O7QHXA
Js530IuA63Bpi5rZjx/bDQqJol1j5uQyXmJxlNE7SypOhnNIwLyNFL3lNZAxOcdhLPgzDE0iVxD9
xcP7FOP35FxUvI2dK2IMm6M5G4I/3sxWnw4magXf+InBwec/4owYiTcVfkeds9f1CUgYJZbfUnnJ
H5Y0AniJLu8Geemu9lUVbC0INuPc2c2fns04HQusmm1ZR+WAA/Nu9SiwFlC/IBOvvvvROu6X5n05
L5lcGo9nsOKAtdz45WTctjl/fvOuW0PPQYhPnzVOufoxXxVn2BERxNZlOLh8akGSA/xNiarQqQMT
1b5i7jN/p9CkRy9U/WqJrOy2x5DAeK8TaTsmI42dx6ONuwm+3TZiHPsyaanCYqE7pMlZcHcjpOJ/
U9EqS2w/tsQ+n9g+DdVUsVLBNiPRPqzOWZlylEJEfsojYU1sm9ml42/CqzToue3m5RDzm2nXbSx5
6zhW6X9MX+SOJpkOmh2D6AAxXR5HDMaipJYHNbE5aLqhQxVFqFtzrcGxylUCNkgJq+Mzd8nzJKne
TED6E+3pPOx/Mgg6MhqKA+BX6XciNwN1bbcvLO5vWpw/jUbV8/YW+U6BLie5fHDE4gDe9dHMs/v8
DI13OiFYpeFEjInwdk+FOVF9rLwO00EXaI7gCmBZWYGT1m71bjtreCPlepR3ryOYeGdcgRVUBQHT
y/Dk6BGb6VsS0XBJRg/mxU6B/5J6MNApztv2syDzd1lTn3BI4c2AfFsJqOoDjHkr0xdHhC57STIV
IavJd9YIUw72Q9H7La6Htu3tMZIjmXTZeWhxzRQwUsMHqhXdHdeUSZfczu36Okr1//GP3F7ZuSWu
7zSBuGgX5XrtVL3Z6xYznUUWXFeqyzd7N5WmnGJ5zc7zZl+eYUpXBZNqfIbGrj1lKSE4d5AjoYbG
J62RgRGO0g49GoAxeZGmqHmGpDTTkaFNd+EH0u3UsShW9hx1nFGRE45rMwttUYGayL6G3jWtjUjV
kquI/APwDpa3GFZmKuVICcQGaITuxYPAdwPB3K2sET7jCSwd9XBLCgT57ZPFslQSVDtEjDzxTNGL
VPzm3tkL/LC6eHCz349sDa/MaCnmhd4GBT5wv9HIBA1V5CRfZxPYswwMTQ2+MAny0PAhDqDie2h6
SseFJQLgAOSftl0sx1D0q9rRbt4u8GZA73eJNbUdp1H+VDu2wjZDrHyrhun3237AXqaXNrdPHIEA
YgKMwkb4k6g7QLjN0IOK/zDysMr/ET2rz0gGYb+5EBHcmvqEEb+84P/cC7iZJ44Pt+uhgqn7qjjX
PCav2++H3Inh11cT3O2aEZDbYIXKQVbZC5zQGeABA+4JadV5G5mlMK4JzFkgp7MZaszwk7Yuc5Rb
Rd3xzcFvka4h+R+tWCQBGMq0NHuLuzVbQH7nfmmumY8/iYmnNlvkMcj6Jrt5oalwaQO9hWNXDDcN
6XKQPobfO4ZJ4cIQ9L1o739KlCdKQLZIhSAqnM2DB7SJw5PQypcWjbYmeJWUdr6iOiv3BKoLHbyX
tym7I51byICw8dgLg6/JqWqGpw0gKIv66Enx82eOH8+khHSJVLzID1wD6z1jFgormNnnEQwIvteO
7uPomX26RnbPNTmEc+/fTBB+n+FScE4Es+c1LA9kyU/VGg+u/LGIhb48rrtAI9RAA8SUL03YCoMA
K/bCSjZs8dkfQ73Mh/Xpl1Gc1f4bjpW11Kej2gx3UpPwzjFR1AN92TgfjAXr3O9Drmet1/XNKdzL
LzbxzmKO4KI8VQP8T3zIELAHkkkqNawicqE44b1UPAEi9Yhvhrd0WREP6gI0asJZs/N1EcgRmCg7
JcHwV9xYiB+XkQSpYORN879IcEHUShM0S+muvfrxgINQfJkFS++5ZlxUq8zZ3G5QWeFb+EKYnGvD
mEm6AYx4hjM6RqJXjVEv9PplxlRkSse1QZ6OItnl71bpD5gZzskZ8gd35i+uVZx7NdhcPBxQaHDh
fGBOOgHrW9/ysvT2Tlog6IikelrGli+sbMlJwfmUp60Qqq5ZOngdH716yIW8iPD5q3ZzeIaBwNXJ
7W0gFXUq01qivUVfMDhZnM/fsfJZVgTKPdX8dYPhj9k+t2zmv+pc1eQTZ74ZhGfFHOlmynbujPtk
np+nCAIGYUJr5ImJoCLo/jH/Bs2Wl8ocM53XfDq8GPBoqIqgTJdKZ0aTvsyORloefBtw1FKwQ4qK
Tw37fOXcoZZq/yx6HHR3Wz+gMRW516hNFOgrApBR3piAiuShA26bs/mJ8AAqyseKs53Q7gHvgtQJ
acrX6hpKXeGduWGDjiZkVoHBhcVkPA5sNkQOHRMdMpihcZnjHs2CiJfQfvSL6UGX0YpleYjfDMjR
nVdu6whrIoqdwmEn+RKpCGUhtxWwfuGslCm1yk05EjTDKI7Ka1pnB/59r6T/Z70ssRhu9zBlLEKX
bedH50mqfDNDBhG88moEqUYZlmArznK4d/3LNw2g/I66e0FOvDhI/i4fqveDCXFYlQn1+uLzK/is
sJJhUpR+ynPH9Rt0W4ZAdLUKIoMVkcEn5W0GdWKJJznFhVqWdd8J0F6x04h0OalcICpwqVBRfpLT
sXyvwetN2+VNZDjF8Sls2+ltjjcn/d+gB4bL9iH+HYvXJXq6QREO1oVGDV4xONKqlN1g1D6yzS1d
wP8mk9MY3/BP2W4lPKx/dUN3iWMezLfCfqCXeXH8Pp0/a1aePe1rKxGjZjnOu+I2SZa0VD6Z1nDy
cE+Li5TE0t2w3VxK7maqP38IC/DqR8mxPVfreh5dnTYQDcMnyakA6T7goyfcixp7TtdaenbUxl3l
6JaRGMCxmwKfMfsa/zGDqLQQg0Q2weW+uicfhvdKBKD4TYeP5+ZSVMB3fax84+/PwYlwCi7Yq6q9
7/ttr4TtI5Sm81gcXyYSu5hXjXCGOH9otiwWVKKjrKtcXPDqbEIFkm1Pxnmx3KeRa4y81pAbKU87
uINai6wkEksqk6O/RoRYXankbyfzaQQc/KDHssEAH8OKTKU4O/za4KVDFAKSBfWEOhLxm01Kxl9S
N9jNrJGhHaVyE2PKORC4VK/trVgUGHUbYw1j9fo/l7YoIFJzszfi7ArM26mUxE8Sq66tR4PDOItt
FGEc9wSLV61YSZ3qZX9UgjdX4FJ95OWR742gzlytoJlouuAS5zp2UR5yQtGLMUNMLjnM0qcrXO6a
tuv4PbBWKViFsvwE3SBhHE6GIgWTXncQQwP3hM+/vMOtqSuvG+xBsLKwc/D2BpVxqs7+FD5zsjWG
oj2Q4TG6GGVKrSN9MPSmsj1/N578Jy/hfMOWM/LDNJJXO7prBbE4b0bC6gguxcmhvcQqOKAt1jKp
WIxnecOcKmG73ONlCF0wNCkdvzTVEAwFdhfGFq3w2e1ZfxpzPgMcpU37cV5BN/+p6ch2vLAEpTQR
KR1IbUsS1L1/XLr44RfbnXvhOamFaQzeLVp1m9IEgZdBtFHIt0xjc9D0FP4mZEF5g1WpyBHcYEOh
ssP9hoHQToCkFlWeJqexoJzlrPF/hS+G4N9I78XqKTavbedIe5dide3td6r863NjTt1USIVcdfl0
itRL5qmo//PwsigGGc8kynJzKMPHRGo9V3BE9Lg7Jxmyf8UNSr+MHcnmDPPSX94SgV3L8A+daW7I
zhcgBOoo7LURZkIC+toxT47zKt1oo0DLbosyMX1Ul/04lzsbkFvYDwaQ0NTMEbeTuABjivi5S1Qu
zMxvjQv1+bNh/YgBbjPENsnqAwOxcEInUgCTIkDb3MC5ED3ZKF6LEpCpciQIEoYLRsIDrpe3Yrib
mowzEZeK9uqMoE2x2UftCZ/sBwkj8BL37nehW9ahkN+NvASZMNdACLcT8xXDz1escGzACOIOorrz
CAtntCafXOW65yV/QfmdJu85NlBKRszdhhUHIHCQn0qcXZ4kVndNs95z2rO91bnP1rWUqxMFGLtp
QGHI08QRROJTsOf+T300pq8RUSiYZcGmcO0lvaqhUlfDMejt2648FyqXJ+33GVJhGZgH3RDSMKqk
sgNW0Dvf0vfIGoIYkZli91TJizdNGvI+v9dlcDMHImDw+PZpDHDAqHOJ7aR7oi0n7xI0Abxm/7VG
B7BCTjnR/cJwqTZkHri/qOO+kAhHZt5rIyLOjAgD9kSljIAuoG2h7sq3ZWKLuwTygus3D+3+9DpA
93BYzDDboBzhGaJXbyA2L3fvS8dhgcbKbeiGVeJS45ZDFMnky5dG4gZQLfy4unnXMOb48MWkhrnz
Ny3bm/5bW+Nz8UhSEEAQjFwiXHNluCxduI2KoQBtY4NS8xURhQszIZ7+7pcz7kUxOSR0bIpEcvkF
oWsdjHFIYYk6BzT3GzYp8tKgzcmtL6k+ClOe8JdUApwPux8NKVmR0oV5PHz/1hjj7d9u52rzLhWo
DUcOqthf8mG+MsOJE9raeDECL/cS8bmSiH9SAcurPuki//hOXoZg3e2H45ppCTK9QBmlJJKDvVoK
qtnlXyLKRmquEN979uAcqTS0R1hJLKmbhEVImZqrENY6IFEGz6kfL/MXoeWPFfRHolTrIhZvOQFg
94Fm/Pp1LntMms6iVE1mSY5Bf9scyUgxacJg4Fk2UDBPSe3KFrlSN3CaK7cFnj6N1xvE1Fp7X3MQ
93LJkXPoJ4dvVcZuuWkXkro9NgAszjznsmQt8BebosvjPosoGuz/0su8ViiHScTcj9xlIe2uOnTf
qJ06GvizYDqyyJa7rwO1J4ChXYJ0pOwz0MQcp6S2EAVFGJ90jyzMKvDs+51XNXQNB2vWzOBnCSS5
1LsFHz1vgxBWjRgmeJehdEbcWE0sgewf8SyJu1695bT+svIUwVP9iik+PKKzH8CQRhZbrG5MdYLd
FSWFJqfRRsxwvEOKUy1sFVBLHvkDuiiMNym4yjwarFItyxYq0ZUcmVnanMbztnOPkt2mLuNevGUh
7swadtg6JaaHjkmafb4YEvjm02TXaXfBLomc3j+d0+B/QzJS0dZXqfQyNt2VlvFYDPuG7S54Q0cW
s/1sgMFtwFPx+9Jrj5Vjmudn5tcmahlU01fQwrPhhVl1CTS5c6X06tmYhIqhTBYfTiwdWNLlLxZa
DntF2Onq5evD1bL86pVbOtMhHd2Nw/aEmcI0U4mSZ+ltmqtf4KwMPaSwEf9bAvcyGKmaoerbW5tJ
awLY59kuXZih5YKbfBiHhRNKmi9jj9RftnGw6ty95VUXgKPOyfUlP4lNBTlsJIXRz2EU3zu6JFJM
YRe8FuS83RxkPgvL4MErV4lMkpWkhraO5a+zaPR2n+DJByGp/GHfY1aR9uD4RAXy+OQCGxtKy2yT
cJBEL/6BHgzZR4cgzPi5cZB8j5YlKOvCgCFAgSA4LsgeLM6kDi0jp2pAPr2CRqlIG3s0VeEDXhSK
nb4eFJ20xWdaC++4807FqK7e235yS2f5qpQA+2zztLxQ2nqY7FGskmcnIOiBgdYVbtOA0n/Bkv52
YcXEuZ7jQSS3S88iSDRK8tMrdmghc7MsDJU7mYvZbi3AHH8ypugkN+AhcLRaM8dEVDXU0MzrgbZe
nc1Gp0SR6yHHxw0OzxOWVPC51fshTc+rP3CXirxrNdSQ81wAT1cCmnfhjg48sx10RM+RGMDXOzMm
29/GNf4A1hVojn3CMNYt4BJTTovJ+tn4B6aCgR8qhPNWmz+ov0vIkhS+w5GNZrRXiiBs5fv+FCjZ
tPXUDu2cBYq6je8C1A6NtVamN2ExGVcg302dCTbsdkAcwvktu3eexLjbu6qLw6oMcC3akMF7Df6U
RqZG27UKZFrrTjH8itZqqFRkiwUWCPXf/SlffLO3gQhZkfDnjJF7BmP04KXNer+9Ie3R5uiVzEwd
hQcK0ft0K3rI0Sg5V9JqoTJs2ovUXUQY31cP8fU1IuKiGWTRpWAWcZuV9ITSre61Wuk87guGZ6+d
tgBdrlf476lPL2DBk4geHW1IFvK8Qha7MOzzVVEoKfIJf7oElnPfUwXg6f8Xi86Tzs64DiN9BkET
HY0lk4CuQi9Y/VrOGSRGv0vjMZhLb7Mfz1V8bk0yOjn1WPBf+0zTIB5n0JdEGHOIpoO1JOjULvT3
3gZp6wC9XkltVacUUR3WX6XSFirTtJLD7XCz5TGsKH46VPffuxKteFLz6WfJpEYfYA9eb9WR2g2t
jtdis1J6wnVt2TTwkZxJqVduDLJa4YjJwiL0hS0t+plPBZiYK5Nubk/Pfn/TsmjaqETPegSd29Db
Y2DYJz7ZTZjC8UzUUbEXACLVRIhIWMM+5d/PJmCMJB/Zw83AU5U8Q6XFRJGdZkU3o9ys82w0ezuC
dxir5QNFdVHXv3FVjxwSeumbTq2d7kplApGAj1Ccr6avsVfZuHQdz9n3nL/9eZM78dfcn6YLzTpF
Nu9B2rWYHruy1KyiMpr/rLVyA4d26IIxqgmR0yLHX+TDe0WusZtIZlm4tnKz9qkdrCNyl9StY0Ep
VefrXKyDWQaV9sPaqA7O7gB5YR6uZ2ihvHvwRXgZqmT+VgQmiEotSooIc/feoKVPGCheXdL2GIGC
4niRKE7hmWg6YZWf4xmhWuexaC0Iw2br1B9MlbdZTblHkfxmJbTKFnoPIk1i4wd1KteN/bB+W72q
ndRKs1/CA/dnr3GPWrxCad2PNxATdP1lapJMR9PtRC3hD6u9etwNYMyU4rAV7mlwZqpzMy7wtVYp
eiIb/xTpilqLqnzdBIFpnpRm1QzTigLiDhbqI6TIRR/4zohE7y4cpAIQ2OsN4nk5OeZD2F1cIcbA
3b/izJI8pyVDLtd2dycGao5StX/y1rutYzGxCog9pTTZUlaazymDyCN3QZHWIUJBSRnirmuW8SFH
KvQndQmc3+FOx8BWimLpM0fHnT6Fy2Toobl3EUzujNBYy5uk/FHRoxx9BeyitiocDPhNcSFn/I+M
eS0EqDiddiWrBEGO0crQilz6QTt/jL2RjL7aBOzyIY4KvTCaFN0ZmBM1t6Lq+NSqcNnVl3aQzkHg
cU97qHBvf9ECwrDvmM8DQ4qWTfCAfyFn9rL2CYlbM6tRCN2R9jn5x3TarfGLzSwth2FpzYCUzC/K
b/4CxKCzVDIa+Kg5w9hmuCn8AGSSlaComNGn0dHdwhlF/lYkmq1BQ8sUAtpJPY8KbKCWMj5ednxQ
+JL402aPlcvAUd3cKpD5OsCGYZlhgbtWM40FpxHNBACNM2ss5uQoR2EAjgxLFUQqnZkQPzZqcMld
s0QoKnGjWLIZgMt7KXVv1M8aeCtyOw/SsgZLZ3rqRsTtBmSf41PF7BZqoTQlVrPb/b5IKdfmM/Xq
PWrpTYEDHtuh0X3UqgqjkL0tqFA6mrBYt+mw/sc1Rn3KlUIz8/ppskTB4vmWXqxsCLcK8fSBn0+Z
rK68AJcnCtKDadqMAeQmE6V9d21yKXboUrS2AQL/DDz/VfvzxpP2Bt3pTczAgdw9zJkxjUBg8xBh
1GKPrFhstWDucPmW2mWS5J5P9aVM9daGW4gi1XPZXiI19vo7EFOhR8pP72UPnyll8CUrLzi1c/P4
gseToaf9edOBN2xcdscq66fWLM75YsBltaMnMVKIXEO4fy4zPUhIiEUb86iliCljXdmmNUrKwysn
4kYruCfX+qeRemWX6vAhvERms3MljkVz0S0gIcTUzQRcxv4Z8WkS9Th+Hfd/x0GX11D2X1zZrlKj
pUTzr9Tr5JAGuuNs+gBT6I0+5COqvnSSII99hCzq4kzcNhRYxHbeXZVYCebVXF002mP3pBEdD8tR
CFw9l5ekOJfP9LAsul6Cc6Hs30aObUzZc4Kki4WddP1xJ5hbPX/xnIm8QzY3j0PdFZ6ORVqQmX82
J6XHpKaMkfNMWatf6PklWwaJIJ1h6IATJNr/2XZL52zC237H7xT8WOqdLtl/fPrCrVXDwBbwq3Dg
/ed7yyZoFhERYAqHAfIswaXT7CwIMJpOqxUCL66+lwnYOYQUTBZKNIsFCBdDObJCdfEz0JMQC589
N/BvEQk2t0Xn+tzq3KheW20oBBMfpb3aMJ07m6cRb/0qKamADrFv0vySyV72nKoYBRn7t29p0E1m
fq//Okl60dfszKLFK7x6BbLHX862YdPUVuUidaeijOdS1pIWWw/KlPWUj+NTSwu4T8psHf/qVm4m
aGFq/gfkyHl30rzkHA+bhIj4jpx3LGgohi6XKGG/KEqAW/agnnhLbA0z3Z9QoKUR4q83m0xd+YzI
Yp9udbAa7CqK9mD5Sq+CLwozsp45SsU5TMVCPT+Of1mwZmhbYi81Xxc1Fx1VEUMYLMM7aTHXBVJU
Qc/mlkwz/i1U0UTwqJCuhYuopTC0B+TMGWodMKKLyQEkcxwC4k1BDqvDC56KilxRkFGD1aMPoyu7
u6SGj31pCTMwtWMOpAnEPFcBG8uUA1jB585tCJSVZw0vMnWLy/lXwJVAvHJEC2XFDF+lB01RyRIc
22ssFNplZT35BiqevatXVlQay7lcUOizgD15EwP7Q9UtN+9hqMzHAwp3DlujdYOuZJfvrzxDsfaK
LJu/aROFBhGoyxx5O7Ay7Cx2HEemBMMY0alyLkib5czuM1zNI/32yteJinbbxddpCRmRmEjW+fZ0
OK3yENeNIqX4q8F742yH07oWVuItrEV7icbiQpeVrKmbtv87VbaDoNdf26SUhjxtwdN0VmVffMbd
V4XAMa47BTgwHgq8t/2aqaSbxVGQTjO61jYu2WBWpbBKTSPvkEnhTGkVtVlBZ4lIB1M0Yh9k7Sko
X1U16MBSPTGqx3hnbhyJUslvE+IbubgNqe8JokvneONr+y9sLgaP42cjJoqdm30aZS5M4kmVqnjy
z6VJ0ocvMlu4ZOdv8rVZ9PpgWcrIVryQWrV4ULm7IFhLq50pE+QAD5ZGyvCuDjQuP6RnjYaqMa2+
0KaBaiSAxBaNEFXKcgRl29yNgncE4olxVI60YoTr3Au6nNZYc+L9dFOkr4FbgPp5myvXxOWMjDuc
3jUpwKbEOztn3A52e8QjVJz1K4qF62VQey8TJNmHOLplwqkORofKCeuIp/qf1TPpkL4FgvQryd93
J+ZLnXGgNI8KVNtS1xXgdtogQvOPAOf2Fu5SiOobr8jHPkJPSHrWu6uYY8JplJSY/HsvrbZ/nsA9
hWMjF8fp0sSc0YSiMUfdROphXK0fdF0x2rRNH9SKIuNu3+YShMloaU/vbYiSI8klV1JsCkjjSCTA
AQJlEZ2AWrpWyjc8dfWV/ts0KmYxgn2rwwfUvnWJgU4SpjmHbjlFhnas5FGYmJ4pV13vh+wdnmF1
mjuC59eXCLRxq9IP8tRfQl0pCBaowwRHxRW7C08ZnmR5s2cMGgCCpww3+ZdOLzaZYt5ZiHgbnU+Y
558BG/RvHp4VoScULdIBVV2ST+wKrXhivw3Bxt9q3wBgtrc5U5gUJCecQxxbsXG9Jdg+cAvAWogi
gTmh75DVOhwXrUtbVhcUzjwj57ogxae4lPy+sOWOuALRfI88ZN7vQJlUByIC/TdzMLUSKC4YOLsf
ByrP7Pfz5L/Rfjtxs/LIXDZpu93P0iD0B3n4UDcYpuxMbYs/Y/hhOUKiwtCosNVkN8SEUr3d8wnG
JGThy/AS7aiZX8eR2GMpRHtr1q8eUBhs9fzieBezF0L7/HBjQhAjvWXPUKRvUFsIoG+7tv6I4KwX
ztBKTxTbH9TAp4RY1/iLINDFY65gStNaD6H5uuBWkRFcn1S84yeKUQTlFhAIh876s8+FigsyRyfH
ML6TTY3RK1dxwRBwGlaRDdKpja3vTEdfXXsXEa1nAdaBCYjtnZWK8FRGguJh5Gtzu5WOMa+PtbsS
yRZPF2vzDg99lSQpxzBV38LYiW+hshpMNQeggqHKltHY0iVd3gU5tbM/5qx6DzSPb7nIFTuyBNLu
VLUzSKPqJHawAzjGDeD1lTqXGfoVPpNVsZyZdtIAa0L+4wcOBMxjQiiAPhoQ7Sk8UtM1o7X1BFZM
UoyiZvXz+cIGBLJ+V4Ra4Iw6ajfMfGSroiZGGusb/HSH0RZ6TQeqHAsrdONki07gNuBniiV82ML6
Ew6X5KXzn3mvyhtaVthTlNxV2gxHYzC3noSa4OK1W0vbuuqFQN9+qxZ98EywFXSUq4LFmUSrj0CR
CvqP8s7iY8GgSy2n8mREhmXrkRMkzdWXSN6yiQsw2bc2gQvhID54xOSV5z3BKVf64N8sVX67x7Si
IBNsbk6pdX36TZk65n2qatXqaEBEh3yddaqrJveoEY95Q6Uc4b6kjr6y0TwiQsTtcvEMNUAsl/Uo
ZzLnL8gEXUhiKc6LTIDsPsQPKDCdo91vhq9e9gUcv4FxwxeUSsQ788S7OO/+60pbyzDhaPn5dWbb
kjtvB/qvHkzT/73sPkgZO+5dmXdswM6AZ8LEEDAlw5b8D08RQJv1Fhvnb0c37l3Tin+eHH4kVtYy
ZVVssCFIOUxtKCP7AxUyRYu/oLN1R9a8kxJyJG+y9HYqUk7cYx5On7QfkukMEKuZ/7iUSO4kdx9T
CixWEaaiavtDynAsoXIP0z3jBoEoKacJz+Ujw+GltMEpXWr9w7ksXSeGyHWdhuimFPkVFaWlT6Wr
kA1nfYJivncPYivGCowQwy+siwb55Il5Ewuee0nDpCAl7+KrZNZYphAU12XG2rAZgeh02g0O9CEm
O1Q9/P8Xab+nMt6Ss65XTtYLHzJ3prDyDILm6ob9+tdLhdUvAUy6xYtSnoQrjYqiynV1ogU0I4Xu
rcKVc404bjy78DnNpeQGCSh3qkFsPFPQ80t5710ZsQtVl/LEOsXop6UXGJNnOqUFKuCcZSTkGRYa
ZeNhNlzpsVbHsAZWvmoQDjvo1TTR5WrrAvc8RvuWJ1maOlLT+uDBKxjzNddUJB53FHhPXnE4TPpB
bBhDpRjWRIuVUZFBUTuxtCtROTme6wibI9sBv0laVJca/3RIJvuBto6oy5xzK4+tdCqPZg3VPhRt
WST2L7oMU8aohbTD6oBEZxgLHn+Z9mEIfMAQyqdQSSGGSIc/lvGUysfKpsXC56GObK6fOJNIll24
SpY8fIqG/sVetDytpHqP7wJg/Kz2E7t/YU5i8N6TRy3G74S7H1EzvLieOXAU87Zy8yYs69HxoTYJ
H5o7MtjbvTA6VHr1Z67Yz7JCuQv5ZX5Ab8/cS1xzaCuzlTmhTzVq+WnQyaCCxp2FHPtFQySI3LiT
Tc5a/JJVYmPiQ8/PIS0jsAMRPGCSNBRlyni/YYB0sGKk8J4GIwwbRXH+deRf7/2yO3KZmU8H6GDb
8Swha12CHWSh3AFWk90A5S5Lt7brMQ7L5UEl+bCGSeyX9OhghbhulBGE6vaATGwSr74sn/+8fEor
7MLNZaDGY6aU5BTwamJGUuGPdk5O0xbOWK4dH18mzI3TCQDG6Wbjsj9a8R7ySLvu/NLSmbjGcIDF
CaX3aJSrfiMuV+n4QGxv9s+Y+Vdust5dNIAbVCCZaX7BmtVGyTkRH9+G73sYX8GmITBBNWObn00p
Feiek0gho49Iewt5jhbWFbqUEugCQ6z9QHITIFRZRBWQOL2yefuJfmmZ2NkdNZRW4QAtwtB3veZ6
t8He3Y6FXv0q1w8nSm9Dtu17njU2T1L6M8mth0UkTe26iO9uhKb/MKWTtdFdpYDBWaOK54/sT0Jw
A2dYfFvoXofLJmo+mZOm4gKp1Gt604dSoQUa3YQGomGw6fYJ5N+lLQAdVnEF2zLEBNXzj3HThp7b
M1NYxy87
`pragma protect end_protected


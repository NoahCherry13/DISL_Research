`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
hvQbM84jMJZCyA6H9U9Xg81ynS5ofGGXwePW87PvY/LJsbyrdnuHXr2HWSEyBlQS1MEjQr5OOoKX
O0FcqsI4u7lpkiBo48q/f9eRwLYce7ejZoIr46z+d7ezBnes9zdyZwAuWEBdeEQmgFaIHvYXqynf
yDjEhsBwVTTgklXBLyoDiEiqMRGEeBoh+pxUN9rfBNKwM1BREUDDe0acShNccw9tj+wZbuyB/T0g
PBTK3cHULmGMpSMiGLSv6jDlp4M55KG9YGUpFbjIfKYPJ5T3JX+hEgGAngV8LvA+Ha6nDcVp4Bbx
QNGGNaL3tmDPxPMfid0pT8rd9zHr5zVBA5KfIA==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
TbjQJVnBf1WnoUfAw4ftQLqn+2K0ytYAsqeQrQtwOy3rWHrz4IYmW/4Fx/oRN2yPlOM2bIOFVjH5
T3qP4pZs7ocNUonD6MygJ5sPslUFza1K5UXmol7RnaPlxPYi+vi+728P1QrXNXN5eK+s99zTWRFh
Z1kepC6vdQutzzUT94AxeFwZF6uV27s2xMOYplFzYUj0GR4XdCw7bm+3mcPIQuFwkHzVVLwioBpU
IPMMiTku77R1xBqny4UDNag+/9424CPtpyeN3iRs2iTNHTo/mOmF8kjy3b0U8Zeq6FnyRJJNmJ/Q
4Mr/rNwIH4mTZLv/BX2K9W0wBWk1LSHr46OqXwAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
LaujgcYJQD6EwtO8iT5sgP4LsdOeSxCX/TEeW0LTfg4NmEOBJv4ivHbe5j4Rps4Lv6oWMDoxRwpX
nLau+f/eVw==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
biV2Sbv7EzxvkoRpMEHGGPYii7pQS4vMv9Mj/WVl76ATNhk+D1Ivc8TtdtWmrnquCA8PK19neci0
IMSJkixt1I7xT/KMNUrAbDhFKJv0PcuaMk5zqOXHmGp+v+a5t6JKREDI1OcqXE4N/O4zp4eg5en0
TjVeclqwmklJAtssFt1UV4utfvZKz7PM6uMdiU2I/G6qSlM+wGlDbr58LxLdliMyMyT+nYqvR6P2
kBSjohRs3suqJgpFtS3U9RsLlzYwyPz5XJOvm2YuDEVU1biW1xFAxUfhQ1YnwhAExdXWzaRoexoX
Yl7A3o394FUyvzAd4lSWXfSOhrdiiN9VaJEjAg==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
lJTs47vENtVGsVXd1Eg7C/TPzf3mnhs8uTayhC00eVFkHp1rC+ltQt4OnOPpCrFWxiMicD1uJRzG
aQb5hjkxV+AbTMb+5EqGs6I6LZnb7shGX2H7Awl26r4CYT4ZIpM+pthrPM1+9pAiRA4CBdhfXuCu
kJKMXx1C9aSfxcp8MghYgPvtm1sR5Wb8FCPk/TRg3tFxbyX4WBrYh3aoHqL9BqYhWJ39cQ2EIA/i
7zIHvtfyiQlHOmrxDr0N5aZ/0xkxiRpZqaeUXhW/f/Oum2qabDYY4fDwbFKmViVxHhCFy5ZMF8F1
dxqux6aW18cCIFWpGnCLBvXg+ovUCFqu9isQDg==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
eV9Nhn5yZvaqBgvV9xw6p7OlWrz9u+8gcOhMo/gL5s/B4BdEmHlAUDk5sVelG8iK7APLuYz24t3B
NO+97eVueLEXJS9eby+Igks1DIEfDDlPB8hioNlqEF4rUFxK8XVnmHublmpHLLfMfzKDbgRcQCJa
d7AuJZulhbMUUDV0KGs=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NfqnvST7Y/WY64Q14j6uiRtD3Iz5cYGv/qlGcERYa3LlftJLqPwgfG9Pl+koYEpsYw+nGZ3vkBG0
tnMSksbsUvghzKnEgv5qcJK+1W5QxDAdAiPzhHDN4/fD9xQjN1ajpRr6JntOetgjkWV4udCBoqnG
2jwtAJ1dS+h9zndE0h67HKWgUxiMpAzJ0NqPt/YXReOM3d/LDIBJHD8YRw/bl0fV3rrMpdXOXrao
YRQRF8NQrHNziSWM5SEKfH4yG8fZVSNNBEa5YMV8JomjL1il46/cf5/byCFNncUUOv0mx1fbWqt0
w59LdfXVwZoxKz1nafUnww/TaxkyPSe+MLkcdA==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WgYvmNGO6B7dy7b+k77YoKoKgXoxKJ+1mNOXX/nvRiamPL3/FHG3ved9DHgmyptvPrSgs7paPQDo
dLyN0dbBqwUEZ/tfeVUnhUNfv1Wi76WuwznT9OlqB5FtG3dN14N5T2UbUVDhanQM0hsSqRw1Tw+o
p76mumAxCZcA60v6THiJIyQiCftAo8civrVu7hNFNsoqrrVJkEY+wyYrxe+APhUb4OU0r9/g2S4Y
O1uWl3SenBsFRP22ohFOIenZ0aU75RRW8Xuvag+q6bn9AaV79Hczy2FdFbwLdReE08brPtIs3ESU
gztUnTdYw6oqGTs/k/7eaqkKMDO+BbGegTq/hA==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ZwUsAhwZiYf4MQzBMVgTf0WMgq6Ejh+45ACqL/ECZTgaz4C8SyFBnSgu4U309pHMVlja8CAjuUft
jeZA7F0F0aSG2+r/utsjS18sfERmIfVvaOVuqJhu6WsfL7YsH5L/3fhbhIGmj00eYt8x3uZy9dkW
lYvprv3SMNp5mZtnfFM=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_01", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SDy3G05ATRMnh67HbPbno9++CDahHj1HO22h5J4Iy6ti5ODju4oLiKfS/AcLB5RklHWVtRBYfeo8
SaGszoCkLwhiCaDTEiuK+PjlY8SKL5Tl6sbrmZeX0S6DwJYLQxLrFtcNdnU6IntTJxSeQk9ADFio
yrmhCMiyoKqLSJ4LAjADrcVRlmuC02WbbqXpLcE64TeIF6ob9azDQhuJf7Rdk6DNz5voC5XoCZhn
niWIFWQWLGjn9EqaRVyCJE2scpfJqKiUFbhSnPV79bIhaVG2vZCANZ8pB6l4cQezvXYDPB5dWzLT
2J1D5GzPgx+Bv17pXTkm6WOihD2N6hB65zpKGA==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20640)
`pragma protect data_block
8KDAx2s3YuYjzrs5G0E1nKpCUMPi2FkTaqK3Zs3tYprwhTJ4Qu19pG6xaWAAmw2S0idFSqCkFOoE
aRA+wermcZ0NbgiHXnjiC4xVD3LGjNnDW9NT6GR6lBBsZoSRWWroR9Sl9Km4JFKWZ1/Z7ckBVNAY
Tf4X2nVNmZ3OCSdIltyid+vlOit3GvodzymPgGmql2rJe1Fy5xHshqgXwCBOTwuM8Rn57qyh33JE
Oaeitp0A7KBDPZ4JvzfpBQHj9krgmIK/q6wHuaISQwnsW4XOoxFJR9bA2fhHhZzvqreFPCbScGTU
MnRQKxdQ6sJNFmaG4jXI8U0fKnGJM3i8w4mRhlWMMW/BZNg1acOaBSrPssygXTOLXM71v/PVDgMJ
CIlWKItauN9tyDloPB+IlbLPKWWALslRYx4BmyvkZYvzabJZh1dmCKwiRhV2fJE52l3HWF1Q7T2B
i9RXEyF4XPH5UOe3CLrhBs/LU/bYLa+s7pWg/jHi7maZzcRBV9wD77BMMsTEU6IZvHlKX30TKSwJ
AdT0XH2eDbmmWotZiYp0wWMp602R2SVOc0j8DtMnyp7R6gbVVehCWnyXmvzWUq6ShQH9PRzFH0KX
ekum6Det9234qjLeMXPKyxe3pHFA37GbSfI6y1QGoed/zzOtYdTh3PGI9yge9wxAPxwfwex70GhW
wG70pc89RyYbYmMmJdGMZb9fbbsKgN6F2A6HgmtocM4kBNoN7+y93asObb8ZXKgJE2SkSLHej8YY
vLwPtdzOgbNmKCFLhoTmkfb22+DlY44Ise/qY8AW5R+Tbu8no3aWyz0TeZ4lmMN6HgtkxG5aX59o
dI3cqmvSMyFiTtY1dQ2D8XraHxTep9TvocbmgvMmMrZGQsrSD/5Bl81dK1cK6stteYsOgQXcnB+v
Ug+QMWazL9i6DL+jYuH32Wv8/huHMyRgY2PI8nYsQSI6nCa5VC89RA6s2cPhV8AU0WrxAdUQ6VqA
WGd9EEd8jG9+zGB0rujPwVEz9UiS8N3FNmxhOyYYiY3QiELNRoCfzq4LB9euajTnXwDouiZVtJOg
mRXOrCJBd8nXwc1vqMLHJS0fjBL5F+efCUC081xYq2g8c2beyf7pjwW2xOn7v/BzdICrpos3uhR4
bkG8J5qQg0oVdCaFAhXbhl7YWtdipuXiWhY0DGDOMK96TZHN0mMrcUbec3prFoziBEXZKe5xsE6g
doizqmBNtazuVgmfhKtmF5v2FyuLCSnrnzyGAn5N4UbMWQ0mUVgr/colDH/VzJzgZKJrDhMI49nz
D52VwyEp+ZUgTXPCwFzPCBwYIBTGTHcVTgMJWhqrFtyz1Yxr/ehBdSsaKIRNsH/z3kuRi7YT4CZT
Yo21KpjWF2Johb8nmPYrv8yrC94/Brz2lRsVugy6BV3FDQSRshZ7qA2JhX+YVLIut4WntD2PcD8L
b90mAXbxNMBnK3gQA6Cl7boPD0Vu44wHwfUtJTS70Lcn0oYlXK225eLnU4wui38ho0HPtRQnCzYK
rd10jZtFIov7sxlG6PPGmUaXH0+L6szZKB2X3Z8iDCttEdGUCiGGiuImhaAvTuRtPzzU8QCfLMK5
tpR5Dggv+K5OONliPmXx+QyYrZtlYkCLJsD8ic05Hod51qCCub9BXYabXZhWkKQZt/FBizz+62CZ
+dXYq1+tkSUEv1pVTSFkno8AwIn/AR9+fBOKIUkj/2wwRWuV/HM3cStlvbrp/tymVwRHFmVHv5wk
k3TyZgXJAiv8cHh/H8MKxKmuu4Y64yOFncFQRFNtJOO2j5qSSu+GPy/ngg4ukKaEOwBwfyH72vAv
NTOxFrOfTyocYAYguw8Iz/bHPUP1QxPomVBV4S0nwQzVW6QIfjNjjKhf8Md/aaJOT5xLyGrBASTZ
k0J3iNHIII7sBWRONiRjsiY4SBzu12UjVGOkrzw5rN0L0W20ISQI4b6llcayzPwvik0QFbqkdyat
v2g8re0wAzc0mXcs81B4j7Dr3FtHMumcvvzIS7sZlQdzKxiUhydyqYnKCGJ08wFs0M5xyLvOtoBz
UFOtebv1iMz4M43Q6pi6i7adb0hQ1479TZ0w1KlSli6wiACdgGOtJXU1QiczJJRiUiTpoY1+3a+0
wZbqHrUaOOrZ9g3pOE9rsB0bRhdn0CrthxPKReiqP2NPC4HWTnQet5VinevClflHi/Jg9NiHFLVk
mFt+UPJgpYrDfUN5RkwinYBEPhvorjbXLiXXKyGphz7xx2zTPuMwiHwWP2JDp+ZIL+juwMj9/rD/
wJpADQkU8BKXsKE6k/fhEDxz5dgJCh5jCSZTwYcjTs5w4brY0S+1pvrd1/JZnEtuG9jdQt0xDpx+
0zs9z/VDHb0cBM9WDCRcCfl+sPlb/ltqHFhsrF8nYzdTxtrneuuTki/Hdh2b1X4SchToVbHm9XRu
q9XEb4Jpb4CLjHDb+aGF+cnbfAaGQu8njjE0AJhaQ2CR1h92AsQM7lpehSc84Rw875pv65uB3NoA
yDZWloQ/bzzimi2L9TLSGpNUwBq/MjmS8MlXv3u4CCvunZQsw77/U42/jw2Au6Hd5JTsnoXkU3ej
4h5VAsQgXrypnyCmwFOtKEe52WwcybCVw01sGplXG3zw2+sWD9UTsDkvqV4xTR+Bq6WSCPDYzK6u
9rZ8aYyV8WhSVwvHfgkQptYjpVBx5Cr3qIgGnFU53hrYHA2/Lkjz3LcAWZUohCBs8h0abinDD2cU
TB8OJcy83Ju+T5dWp9k1snockN3Bc9PYxvmshbQ8L6ViFydUyfs2lnHYxvCaNnH8v/YWu6QU9DHk
qTTnNMQM82Tekut1VlSb4Z2hKun2wirtCL9eTWb0Qs0RoiR0HJTthO44xYyfU1a9HgnYGHl7QUqm
2bCgJUogUfGEH8/XxsfKEa7gV/q5IwGRxcceFeey0/KXmKHVvHeKSrFBf4Ugn8el124muxbOHGxL
6Y5YUYAWr0fAyO9l11f7Xd+7Ln0CTl2Wy8bGkUc31mcB4pMwBMCQYGyEeOyjwfTxwPwMyX89N0tL
1ioJFVtQNS/kpYbs09UlxK1lL0IGoy15O9zNmoUadbDyqNlXScWmIVwBfViGz12F+IteCm4A0Xuh
7BuRaQimnEUSm0ziTVXRxrET1sK7E3kNBgpbQPP5Tip9V/RiyfFaPlEPWtfkrJzpWk8HNm8Wox3C
wr/wAnUg18iwO14NpgWWgRTT7qo5PTztD+txoLQJSplt7c+EK0AIfwXG5jXx4/2eGENeqlYqQmXE
QOQz2VRSgllF5m7ye/1rxRDvM7kxPs34UOqGrGa63cqYpG/aCNSjcoBSuyp+8xhYbFGS0EAHB2xw
5nEHn4ESKoO1v7L5jvXK8L02bg/pahqXmAdlc9y7WcClmNs2SnGb+Fy+k0GBmpmhcyZ5A7L37j0A
1w1raxeOzQwyYY+R6wDKM11FoJo69tG7DdgT9TQvleob0XS+EPc7G0bPl0IaPtxm5db9MSNTWma8
+xcUAjwDlVALnJhozxxW2qlJo6hrNmcrZY5Me2EQKiPrjeg5fLGvFgM/d19gPLBKfVOLkO0jad+g
NTcNOEjJP3BMluVmUlAH/82rnv0iANUBb8W+s0nL1Lo3o+WD7eCEVQnmtOi2DSqqHA7B8Ru8F569
YDD8sapO0MbWPgJbzY+SB7n1qMsuN8QIQ8j1P9NQTHYvnCa5o56p44Q04zeic5ERcq89Ls0S/i9o
Liy5YdWGcB6su8XDAc3bMMqBVX/Vtu89po1AKy2HlywU/XOMTFk79kiB3m1QmPD8KOmaAibcuvSy
a4Xth4mct0fUIiNUuLxBMLt5g6P6C4XvbobMMLrKTPc4Jd2Kg/UXo47kM7Fsj006RgGhzpVscVS7
Jr+oT4/HsMzQJIY228poz0m2outARP2VJI5fHFwuPEA+WBsQpWXjYU2+6aAwakOSFnO07uZTJFw3
3vCIHzIcgsMprqVeZfJwNbSkt1U4l5tboD94U3U1GiQ1JwR97LOeoFv5ywVCQMYbUgQxtzz5sG5o
8ab/rQTOTywvMUw1ndvGhtH6lvwQqiWgILrs/TpOYgizRZJ0ETO4mgXQx486JkvjXoRiXZs69q5F
AqEk2z6RlwXs5RcHFbcTREJU2wRt7w2Evxni0Y5jYeJdCghRwg695Alk7gpuqzR9bfsOFhUYVdYF
RMBMMjemoFcuNkDkI5buPms649p9QrLb97Co4si/HjccBzpdNbK/T+4pW82dPVwQq6aAr7Epfs9E
hVq+QDCF3SDd62iNfyL4iTqK8ntouME2nOL4fbEy5TNGXulyrHltmCuhYtQRHJsL+kUQzOzEyICg
uPXBafr8Ke0+n6CVAtlF1h1uXa0wvxmDOgK2eT/iuc+emOhiuDoWM9z6RmRvYuBYtlcwu4OCiG3f
s9zqCMbQQendAey5Y0IlIBqc7yDDROcOxEP2Xdm5nAqNDNpaDt6gKQQk+V04Jq6oLTtiERXiOUj/
zKCTRSdkz8ZYUroxASx/nqrNrqWyEeGnCSG7gOK5GnfopLguepC40Nv0aQ1R1K9l4oTucajlognM
gV5/c0OwA54CtKpgdSjh4rackm/kCGC1ql8HbUwMd5yDR6G+6y+JyEQcmOhBRRIvw0imx3qfsTf5
RTex0zsV92aOt3QPtAPGcKsdfmWAyteOQ/h9r/UsGz1ZOfHgT2lIOwRwaO8/pi/xacKQ22nvyzk/
sRlYAyyiYI6sGehFfpD+6KLMXo8ZTFHhzOtV5ArxQYd377Iw4OkAWJEgVFZD5VO0youQ2HiU5z4v
BBn53EQHMeD+qRkrwERW/IfdYG6UWq6Jm1U8cvW1od6LVoBiTB5lUCNdiB2adrQk+mXp8do42nOJ
l/Uua0qSlUbW7wCD+x2ou9CPAWTjiRpSNGz5Qc5nwMo7V0rca/PKHMaJYC0sadVTYpkJR+PtKE4i
EIKiqpxBCYJgdMZKVngND+kLipT+gAZFsXj89Nh3YgeU1Mjo2FK/FnmZ7SHTGFwWgwQIDxRAxutO
BAKMS2X/0CcP7Wgb4M8ubFt59rRloR3UKI0eLiIMjREPes7Vexz2TjN3m4u3w3ke/xIjlG3o0t86
gvkXuh9WCraJhQiC7aWYMfTqjAsXmdSDqZs5Me8YRGi+RoHRUypKiALxsKIDkZF3DWrUds5Myblj
yY9IbLOdpwR2LDF2opu3MQfT5m4tfNaevra0YO3z9RJsg38sK7oNzWnsqdLT5cY9nYgYERodoFw/
HFlKzFlFegxlUOrGGmr+lj+ojXmdsQ85L7h7wvZF+OMdcEd5oLueTDQn/lZTpt2G9ZozMudWIAKO
QxHV86RBtSSNufPDN3M77Pca20o8Hc1L0Zn7DmMhWEEbERXvftbB/4b6Dl94hgzyTAa3A0xzUTW8
sLbn1cDsVq8Ac5cL6a+4ky2F+rTAYNDSURJ7lJyL7M4q/dU+Yi+3VxFDsL828ztvIM5Jo3nyst6n
NkX6zLbZ8IzXX/2PqRAlzgf8VVVY1xMt9Ar3U1W7uhXnCj4HvX8QrHzl+vYUGvzXyNjly0fG66+C
zfYZ8hNbk/pT5RRoIPwQSkP5I9hT2fL0104MKBHBDIfkKOHCRZQL8tlN9Is/wsowoG4F2hd+5xe2
eoi1LuxrRlbKOfYWZwVWc2zgra8UG4Lwfp63pOrEmxcaUTWTgbkNMloxDXTj7r5Z/a3uBIipC9eL
wydE3lAGKixwzCjbvxcWXlcBPOZQff65CVsI/sVpmV8NnNQ85nWLrmrkbTD5/58tdqTXOpQVLap1
zx34CSJC6UUwwuxv48zBIcoTDfJgg6O9VCxPYk2vKyfvmTXgL0TV9I8dExt4SsnGDJr0vAh7nMOT
5K7cVJVpYANn4PK1+fOCyTW5MsqLVXAWZqVk+x3N++S5np+yiz8Im9ryrd0DP6yaeXqZ4fAheDSz
tdoyi9QcvHW468nk+TD9lu/uX9f8yn3Lmd3T3xjR+vM/Fet/2Gv8otOR4gArVrIvjIQr58Zyh7yu
86wgPImyh0GLcK6dWaX1JQJ7T7ItlUbbZZXFE5wpnsYNgfgwzqj25dVO3TtfiuryDu/OCqBWuUTe
gEczH4NsrMtJP/lUWohDUr7FPQ4wcuZQ3iv95kMJqnCioU7G5JiiFeDM5e/kCNu8n4S4ZQSsYru/
pFEGaYIYomyBUgiTPOn1z5PN4KsPtn+mxhF78mBhMXdFkGKfkpfTYSpyM6TUhsR/bUzHbeEWDKEY
nQHcPDPivLKRhSou8yfWXxTFJTQ+ae0LaNEaG1xpu9Rw2TPvZRgXdVwfmYcE3lHi/3bE5JkYdYnS
to0PaZom4LuTv9tiEddo6cFypfpdyKki3XP4hNoGXr+XkF1d5UXpHFCE+5P0UlIsFvGbuY5SY794
zc51FZzi9d1T4uAq7G745G65b1uvf39eqEDIk3oe12tWwrKD8LeKQK6wKbjQfmmza4vgb/B4+C0d
iq82RzHhJIgSZAjopEX4nd9cF/YikaPZ/38+w5wTL8nvOXyTdGjmeaOvJphwN2DJXIT/rOeSTrG+
sXmIgV3ak0x5+QImfdLDY+wEvgFfh8F/fAKUBazlAndX6ehhbmjxDWgML4aVnosA+poE3nA6v5o0
olfg8vwnRAXKnNVOtZ36GQS4cxz0+AzmkiFLOdGTNIgx1ArudfeIG8KBHMF2jLx+gEtKDgtaeHCD
ZuERj/JI/BTrE+FerYA/LrHI8m1vZeQ16m6EHDR/4Hs4TUn/qv+vGIK0Ur4ygPwLvexgJmAy81s/
BW+vi/YCUHXbV5G8ORUGr4dNjNtAz6GPZB2f9/Uf2dXBH1zI88lZoZ/A9x9AJNWWUcGRotXjksP4
71ndv2hrQ3khtSf6QhoDL53nC/PtPSNBEUE2igArbaNSs5uw+lvUmAa3Rr35C1APZ2Tu16wznL42
x2Nr5Suu2cv2qx4cVeWMODL/DS1vZK/EKoywrglUbbyWr5bpYqcvaVUnmeQhB0cd6KeLffVxN8MY
oZiyA892E9V7STF/TgJkV0uh6O8X58jkWpAY4hu6dIUMnuFVnv3R65Pd89MojSbSif7PWSQgsqZM
ZmpPq2t8pWzSRogDsXc1yh7MFunmjdQABiD3dPt3i+viNQglWCqAOaYEkp67s77xeWIPpW50j/pN
LodyAWQuq2gVvWbtnIr367wfCfdLtA9iyEsu771KXtSuseX0wn0xts9nlFKZRqiz0JoM+OvXyrb7
GLpSsTHMUrqf+vgGvS4BlfgjZqZU39LwNo4wFXPGN/RyMEsguzI88l4vahWgxmzofcTgIDwO5LFU
1BHrGUTLRiXHq4i/XW1hD9hA+hsi9Lv/XyIBOBwteuGuXevMI5wkCtEfh46/mi5WN0DXc/iTrGsm
SJsE4MgKKQX92o1Drf++6ew+CIwKW3LJ0/JtYvJdqzk84lQWUvezf/2LDWRL7Krrhw2Gd/CBbM++
7DAN2gJK0K5I8Chqax5H0bJ2XekMYWODEtY+qZ4xdTQfdCFMvrNKEmZKLMmuqOcBvcew42vm+YSi
F7t4E1gPHHCwU7gCOT4Qz5VCQr+o6kYr+JauT+573cyDWiMmazeruxL9ecUxHveEKABnyGR02r9C
G9SHBJKDmL3GocGdb/B+kcqEJq71nPTzXemWnLZBuPEKsNftU5/hXZr2BqemhQalH/oehnSeSRRy
12CJ1PjB2dioer0DNjXWF5oUMt/+n/fwq+STNUQM00XzIkVkFfBYqI7821MsX4oqgOPAxpxyOt8a
Gsm0h5pmi09q+Kle+FQLmphdV8TFx3Gy81T094uX5pJYRerFREcsLmBWKmjfoBJT1hORlnK+C8Aa
/3Do2vxJU0UleJ7GxrnOhBugcnZlmKxpTbrhsaPXVW3YiXh6qzEYZpqlJ/aNrtXNBWMRoX16+Iir
pSHUsQkgGNXGJmNtyyTe4OJYpbuynrh4a1bhcO1C739ZSzF9V72MT9lbwjUYE/ozNzWDYsBXfCSK
6uV4CVEIRTOsJRLugvsvz8p1DsU8YHwDno2rTduF6fFFBkiPhTTjno5OaNjKDaxL8dLiRcpx9WZw
8AslPFy898Dr/TeJTTWUewr3ds0a7hpJeTNT3FoYY1fk120GWTAMx1nNK9xAdEvydWmsxQCskhdg
ycFgGtDX+6OwDjQlE76M0Z0ykvbtAe6fqTNxiZ/aVsR9nQ16ZkGc8m5jWHfqQta9n0N58QF+27GK
MWHzGW/FaWx81M7oa/QEHnsy/tILtGIE4FJ6uZaKefEnbsuXcr0N4pZ+f7hd3R7OsJdLnU5YF9r8
GrcBBuWn8OBvgHZJRgS7DNerXlAQN5zLQlo+dhJjmBNmspp5IzBlv6Mv1TpsZDCTFcAuUBsQHCvz
ytekLMF6bulLgfqVqKTg/1gw67Pjkb1417tqOQyOxptoltMqMz1DLOhKIYJiFfXOPlopVzJr09jO
OQBauKoDClvdh+hdD08sFOLazhAyK+JXgDRJ3r5ib5x6OzYRWH27M95lcXD29yq1g9KSsDwd2pJM
6xN+EWIifSdJfli267SmCJv5Xo2gvPe3AlCya0BO/9d9ixbh9eap7dEWuHjbHgeByVE5X1SQPLom
GaQgK18oo7wdDxsvUWFB/xsfTppo4kDCI+8j30cOUhqTMhEUmjLy+HnekKUVV47JoGbECnbusRKn
XVhJCq2+P/QC0KK7veGLHL3UPfDfcIOKp3MJHTP036EOVo9kiotBzShi7iCsQPdtlebI3WeXIlOq
hCBshTw35wtiPa/4LHkyJMww9QohI1tElzVPsIc9SEoGQgbMfiUC/vaZSW4/dqJ3HOlUXPYsbpAA
292XnOqvIuDmIwOBNITlF8dRljLytBmCQdy42Fdydtg/tGheR8clSaJN8heijw9x0xExVl5UxgwD
2Wz+pO8R/MkyhcBWq1dO4daJRRWPwhhpGlC58GHjkAwtw3EPweNXviCW7gbHpLBFHpulIU5i2SBB
baRGfqV9YVsqIpxXOUcvAvtQDye/s18kfyX6bAXrgfKHsppNxBei6vqJDectwvF8hrdQ0dcpik/o
GnQGrBjsrKEmYnjzJ46SWdDP3Dmq8Fgph3YtjrYgrujxNyKDzUS4gACciJJTgjSB5rQ907b5otLt
4Ycd6ZW9EreeKmBwgouWsNXwxgdVRJGylgdHasId1AJG2Vzc0xPBjm22DYDC95XVMv0cWaSOYrv4
CsAntTxVJWprr7bgLM9B9nDIZqErdK1vvY0ESYjhmk3Y6U/oV3COHZfif0ebf7ovC76zQGe5bdpD
/tIAC6DsgDHo6iPw56mltQEjrpryhLUBZhdBl6ptl0GzRcEOcriwTLw0IL2dbDBmqPEgrtBuxjYJ
ag+MEFyvZwQPdncGS3Fu+z+ZF2AF+cv0JXbgKUpcNsmP5wGb5wCZYfo7X5UEmsaAfs/U+HAdakJy
ZZoANYkcseW6iKYl7IROhtuyPAuK0TLmWPZlvkOiRs9Hhc+G2p2EEkUm6+wlihMAPMYwk7CdJHdG
caDBedWJbtRgpJh/25Sm7qitvSqJ/CDfEskdk/XY121TgAlXk9uJ7wqb0JoecEs/3yEfqh5+HfoL
aEXPa6uEGOiOEIQdLcPUpLNbPXYHU6CiYv6S0s2WvQs1MvT8MB/Ww1FHGXlknmFNiONN5SA03zdJ
TIEOxFbELK3rxf8rMAvY42z+E/82Ia3pC23M2eIwTHIJnC4yTU9HE+ev1w9o3E5rfDEinqZXnVSO
jpySxLX7sdtwqhyY7EHP5ZyiLn3b6tyEDm25/EbmaoLsV7z3zuM1C7QXVNnub67mLS8xKP1qakye
nZokOXktnY67qROc5QMQsu9nb+YCWJP1YG+mAwR7Lbv9dpqgGLvFG1umzVwLn7VT7u0MTnake9P5
BwAdfOWmj7XxBsiEMcUNT/GeO7YrVbUElYRtnC5/1BvMR7K6BqYmnysdOq/6bV7xSfNZFBtHowG0
bP1rnhh3XcHuuHkOPM98Xa0ZC7zYlrMX2hv1iK85/m0NhHv6LNnhp39ZTcWYEmr1cqpredG3p7zr
AaOsugH9uZJvts0vBvqLcZdkcwv83D2AclaN/q5YyImMGtkSIfkXSPinyh4ndlLhjq9yyQF9DYdh
ppXERdStG5wWcs4NqKo0F84G0LANO/gQzAvSRV0IWAEDenklkhnWjDHzdC2FGRvOXVnFaHcxHGIw
ztPVOdOTfvt+BakZwtooWw5EL/jciAnGm/iY+S+tRtaK13KQh0h+9sfrmgWL+dBtA/++ZNQq3Ewg
cdijCLRh1Cgb4Q6vzh3FWZ9h+9A6BDx/OoM5UzxC57cAzKzdT0/ty5qUsSjIsgFk9kftkUz61wAa
fP//79IscqM6GGxDaFHEZ0+LKtCXk/2CUyyhXbxfW95h9YH9HhAbfS77YN6mUXxBb+rT76WZKJ4l
WE7ybqeyPWwi9ZpDPXIUwAnDev6LNqqT2hp6fGaTSkDQjkfKBjIKuYAl+4Ly6HibMB8fw3d/J/o0
s3VjMCYwGM9dH4Ss7u2WdMCmiM++dPXTn7dQ4pSgtXrkej2CdTX7LnBQ4HCLAnLiTPyDHft3unwx
hhR94RUwQxcVASEYZAJNBT1R/3Ja2e1jhgLqZa8Vc3cC/LNHF0vMAQ+UOxesv/jPLPGiXCii3u/N
nuLfo9jgQ/uUJnLIDMLgVPKvansPH/7md618WjdqzP+1T6KY+Tlm4AM0LbpvbrnAHVdEayi/109e
46SALK9w9uQ4Mf1P0LI3BlkN3tKz7iJD1uae6ld84uhMHe8NN0/jfeNS+TRO4LnOke3sdyJaUg/0
hzVSNusNmsfQznGPQCOD4eQkxlYitWq1nPujkQQYREsMhgnf4LVACRRsv4+dvtmMNvFGuRNA51Al
m64FcMlJMUFfG+OUtwZpLiqD4WuxRlI4NOVzwbkgYZ/56Pa9Hbz//kk+Zv6HyLMVbtIx1c+b1f67
Od7MY+oh3FWCM8tFjBmr7xFac6Sd/hD45yKf25zzqkzV7EgFSIGtXFYubx4hXlAYeDS9bSIaJZQ9
KFQFBDdFoGx/TlzuCI+eQ4e6xeu3b9f1jbsvQLnK/WJUoqHuZUWLhstwt44iWd/DGfnSsZ+YfmLl
Yy3+qE+QUadtgk4olp558tq386xZ46XNyP/uMRkBwQC9jzbIdWp7WcnyiiX94sEUN1Wdev4WJ7fk
/TFzKJiGVpwupaTO0uVIIBJNgH2eCak0fiFaS736LrJtZRVa3gd/fYNhPc+yUgB7R72VOxnpbix2
IKHiGUwBEFvXlLtDUzypjbwgx6OycAjj21mO5p0JKk3rrzV0xMRBPTt55ztegs7Wl19PPljVdmJ6
XPpvcglD6qTjYk6bQXqGRFxzQnjSvSBs2jitzIxOw6cePjHsw7k3xSPf0NDZmvMUsWxFXnher2rb
K9acq85x+OEBsecWkF5a2n/iwPY636R1q8dl2LuKM0agO1Al3E9j1NSKp7eLe+DOpLSxiKJHTrDv
dCIO9q+/V0fcjg4BlbFhr3+A3vAIpjGtx5u44CCmMLaQBVkqkHCrtJwdOm+4mbEgOu6q6iQe+AwO
ZG8KIaBZaEPVawpa2M/f8Zx9mkCPB/QLVirR/trnsy5Sge4O6xnvSODQSQEhfgWqy9+Td6CKi37V
4C5OgVpbpuwDYpoTxxkyCbHf8uMuWNHOalHq3HXe1vAI+xQoC6/fNiDU6DuPUZWFMSyYetA9LQYm
ZyMMnnrxv/txrpLRtvZPW4BA5YlsOSsyqlK67qoJs/80b6MpYkJdqqAsOgsSobqHwXkZ//EGfMYB
9p6txU0NEjFnvbBfho9w05CRbbp+EvSyzPmEF1GIETtCWq3+fOXIeen7e3xDlGKGOfS2w8rgWNF2
quuUn1YU/Ys+hbxzZPQN/xOuRS6m8qESGejkPebxf5EG8vWRhM5EeFvJZSAe+gSVH1nv7bapp7UQ
AyjHs6loBfXmssxHl9mCTNpq1zN6mg3dOZge2xJm5YD0rwS9B9YCRg0vxW41VgfqcEmkyHfbBU81
Fz9BJJeY+WQY47isxkko447THj6IrpBmFBM9AttesMAz+rwWkPqWbFymUBv7boW6c64uGX6PFHg9
tv8Me55PKafXrMmcth+q2glTV9AFNwgUS7rSQCUto4mFu5sLlCFFky+pMdxHMGKUOUFSokGdy18L
zKOxAqDZHJVre1blnkqz5kxTmUIjTbAfeMxb4bor6787R5ff2BT0x2N9hC63zp1bC8suptQmNtZ6
WHxBTsMhSx5ANc4uWmyqE21Mo5+BczOZW0IxNayWcRWI+3gdEO+IIX17I7NW1VGfiVYpP/bccmRh
+tLVGpCQBuAqJk9OcLcTLb9GscegQ0V+Rh1X41JLppxCpSgxIQFt6RNtdekSZDPzdy0xObKTniVq
dH+PaOSKtBJAhGX4S7hR2tumHeLzcSzOmuLN36euoXyeE+Rrj8PyC2a1hCMn890Gu5SoWc0ZyjNp
Eh97zeqa7Hbo8MrSB6T4iSxfLitE0lMPFCvGP2OxUGMcDHhHRQbCJnadMITTcA5/39XhVTKVFiWe
v1Y4En2KutlfZEQbCLtYy5VGKwWIStUrp6kGFVTtRpY9Tn4P9nlclwnzR8P4yPMUwOBvGOfNwcVK
mC9/BTPTt18m1BFY8jf5DLsPo5jkvGgb0fTku2V/mXYbWbHkmFtr9XheJa9pF6GBtclfQHK0D0Xq
qj+Rtfg8z8KV+kOk53PmpOW4hJUHak9IIbogobvTdITYrK6lwfhHP1I0iCPsdOaRl7klLhDv9f2T
UQImeWOQZbpGq8itlTcwR+6ZZynpz58/Ubu8PO9sznT5VDoNaexQXVkzgxHjpVGyKFYzrtqF42Qz
zD1a0kNmddGNey3d2j25ywNHj0gCmal8ZBJKLWdmGMcXvhb/2iLL7ecTvH5BX6dNJkltwljbIE8F
Fwdox0VxvoBr/AJx/CYvh27Wa5VoQAZelp2lMmFAn+YRu7iNZDRIc4+akrKWoVexl27LOfvEcdqv
fxRSNPd055uu0j+iIZhX0tWWxTHOoiuBcRhH0oXzOVovA0bdoj2HSB4pOwQM/fu/AZIpp+ba3JuC
M5ZmppSgYpi+/LP8cZKMYvAllEf3UuwH/kcQHa23ADfdNMBtIx4wTDFwx+y03HK8huaZ4nT3ZMpd
P8JAFVbUnD5GEuFcFq/sJLmrxQQOAeQyJhdcSG6tFauYfLpF04pmRhrJJQKb/ysKS/Rp2sI4jP8Q
WimY3M0FAuWhNxTV7IkFAxHwK2+rw5sz8dfpZoVQkP8M90c9pHoctDRS0VrsZpBTuydqgVyvYw8g
Yh89G4V7byXgQLHELrce54zMjT1NqiMKzZywUeCcjSgGPNAvyf9r1oOYr/BWBKJYND0zy7Pwolsw
oHHLq9ENGZpeoZeHd7uwOUnY2g+9hQvpe7cAJhXexROb+bCWyWPmcYp6UUddK1nremOVP0TW0FIM
OSgGJcaN1D/WiJwxkt9vCjekBBzcZafTUjtw3iQwsNmls18XdJ9b/Vk+eXg7NpQcQWfeKHw0jrPn
/wIp0/zTrx2TYkE/1QoFqO9W9ELoEIk84Wy4yc/CCL0BgUIs+sKnUMuebpplBNzBE4Yd+mUeteTN
ayrXMJmk4ZIayO11Kf3nJKniCNIb/Oe8Wicx86KO1IhWbVCighmscsAv7C9zNrM8i4BvKWAnht9d
bSQwzC85BZFz0C2zjmwucjKIctd7CMLXZ2pfPZMqvmz0Gp5pxUCQYogquf9YyWc5/GWf0/YXs8bT
l8hZ/rpcP3AmgG83FDrNQDmVR01CTbfz0GARkZCdZfjRzjN7niy0K/+5WkkjWRNP3J45V/36zfiB
jOY7rsnTXpDQVBWIjosQLLubYeOl4Ql63WcxrM8EKjpG8t3GsVj3BNvOKKQAUpMkMVgbl9TZqiKz
JMW1PUF7fOldo1Xm+RfGp7fTCsvl3gVTK3kVcXr+ziQABspX9Rtvv8sii4GZFAGDxSYS8u8e1ShA
ww1gCAxWqy2QkEtH1q6MAOlcf79q5gWi/btzdf7NEQADuFAQQdL/Xb/g6jInnHWcmhFi/5xlQjTF
tIUxZIg4ntWHqv0TNUOOM1YMpCpZQ5lO9Jap/LpUKc8YKml8rWHzdwQ9YSGoCH3RzBH+AIIdmTH6
P1iS3R9hCP7vkLXvtyDMHAVpyZpzVQBTzerwJ/R0TAQUabft1aTBtWoU8SpE4TPbhU54kcN0JEi5
LuYJTpd11FpH44YuOgtRk7fG0Lele/DfRDipatmwbbwgQcPZPt8BJGyXrasSeyFPiya8k46cEv6K
F3nxEIJvW0I4egHFEUvrz5bNVszn04D4JKqJp8A1JLMg4MJk82woHoTAzYkFjLg4ed4vEoafXbVN
Z1Vss9Kf3SbpkFZzNljNWKkVMriOwdNWyFutw+zQpmJeJEoFeoVpdvbXXsUF6CaYYwh3NF7Bi656
0srZpbqxo+cRzfy6WUI9wjLyunxDmB+g2gTvCIDBSJxtaVQDPnX/BZIgsBFI3rbv2F489UxSgLsg
sWSQqMO5YcqugQN7VfiKyDF0G7dOHYWIWzMy4AN2qGDYDubayaHdk1hExXFiFhwN6zr6vfCJUiKM
e16d+vdPp4vPlYlQt8eNRLVZZBFzOCvOb3oE+iqc3Sr1THzviMV26hK21viZmrPnvuXVrgoNd6PK
U6LdgmgFDCkgCrmidrOYhyhjqED7R2qL8lBs07Irlnf2i/mn6h7tm2cxkal0cL2/Se01XfI7PFrQ
rMAutdIfmcVTm12HzoHkftBf/pjy24nmYDDJXgysZhnbIvC4OMnKGr9JYP727bsuvlbcIN30wVZZ
89aQosiBegf4lyNBabtc+TXP5VhpQR/6otGDjtG3QbAtsVMWdAqyp3n2fs1NV8c4p+iskKpNicFC
CVal1MEaoW9na9nDFRCVsmIw7/HbxB0n1i7BEMXOfxB5jlk58otf7wb8QJdgalD4wYGKfZQPOlp4
t0pA0juCe3pDDXqfWi+28T0qnzIo97nc66PkluCGBNR8AshQO4XKiX8e/wuHKAJQGkx0aOnPuuZt
YM53mttiklZwafJ0lJgDtowJh7wZ09xHjyvZddiiYrORSzF1lb48QFlrwPtJINZd4Yq1ZzxSqwbI
VdJLF+Xt9FbWy5/35KWNSQtsMqIbRCBA1F/9lLbiTeE5CLsCHEdxa6n3A+fFjVwzzgaBjR4G16nv
5GxQr0pF9EM0xQ8pSxLrEcLHHmJwHIydHbAAN5HgvgLPtt4vN8OhdfPj59tY/RZ0JGXvWFRXoU4W
E4fU2Gj5+ifbIO6mxRl+YwgEztcSWYmSJhudrbq8V/sWjRJz/0F04BtxDF7GrSSVFjUS6YrpzfFi
6DHO7Ue5sNHlyv8V2rjMLAaTjzbXKAvodp4If6hXSTd6B950Tdox2+jr+OBhRAGnjBGa3gewTXzD
hAmq5Vu5iRqPNe0SCFhohM9A6awI8kiw1q72GOtkxWbr8N2HJabkvcIFTBISWp8MIQTP5ngQAW9M
0xkIX184+L4zwLW8GulSqPeosU1q9jr3r9uKkgv8NZZhDcEaQkSW7925Nr8KRtwjEn6p8TianYL9
L5CVpGe/1N6JB69N4sOktglW8Oj13fcbxeYB8j3432P/xMnOoZvL5Ec38h0y/uY7w4o54uSsAmYi
R764B00KjUoGmL/qGK7HknSy57R0zH7jIrazoCLtGJaPMR3K0/mhdOSOgDI00vxJuhFFmt8tdY2Z
Aa9qlFPA66wh14qCaPItQHfiC+S9FfIrenqwfjTxlgwxfN833WXtSSgV+VCxBdcWSYMT58YOb+tC
+eyT8a70chaCZr5wJ21OBxnS3uGVQjRnRXWebMOghI0KNAE2FIUu1OXUYmN/Tq6dlVoZyNNkJ1h1
1lnslkgI1qGny0nkyV/66eInuT+AncsErHKOT5eA4u3LLXgnX2rGQA+ITRtrbQdzA/5jevSMwWKw
+6/D4rwHPJcdkE9eF5Wf6xvlmCHfTPuVfLWh6zS3VJETtxkax6EpgmOFwUET5wPpGKvCCHZeKXVu
vzsLQpz0JYrYC5cs/gwRKewhJ2O78ii54TjNkc10s59YVN6GWXguNbjmekV49sMhRYtxzGNLJE1V
tUmvusDnYYrR6SuuwWlBXP6iIv9fK5DYrPCgsENoYeLiTUM2gMWjTSrVkFA4NtSIqSIOI2DhhfDN
NMvPSIT1EdVuo2O04QlTyQc8XGI8Wu0VXCZ+fkynivM0XGo5/Y2SF1W3R7Z++lOT4cWs45gvsVrc
KC5Fq+7fauRXY61IWhRgppaXNiwaU0rALb7BS8wxF9sEwH+T/hEsjKFRE2T92yNHXrekasSHsOAx
NiVw38B74GobUCb+HwSVEKBCppxhBbm1SRWS0bSx4L7EtGm+TsK4ylOrE9ydk0pvRLf1w0DC8+ys
Hg78SBiosNf6tAJWWtperCTT4sAiPzLPs/taChwCfqELv3SkfBvjod54ItgfyyQ14HGiuMSndfwu
ZuG0evxBMvc0gB6b6KV4x1vXvp++m+t/IdvWdQoGobVMB9oE+qN5tjfpQwoKWTvkDFY9rVsCbs3V
3eVnlXJG2V6sa0YMK80LeZmd51Ayf4DQUniH6tKPZ5i2J8OIR8h4gotj3Gc/rAWAzrJ96zvsnUtO
W5lkpl7NEmIzGcT01PqfIBbFcXBMVKc17xkbIwpw+FuoCKSKEs/IZTzBdf9qJ+ucsliIqlEKXLPm
wQIkiDVgRIwwaFooUaK6snMj32D58ffmliK6VeT6paOG9Knt43H04TLDaRfeoP7wKvIU77jssGtT
WHARnGNQ+wYeNTsoIWzKze3new8xXGuUxgB+C7gHIkEdtztC7btFih8z1rvwMGpBZ7in3cAeWNvF
N0Ejcw+kelups9IhfzXaELABLdlYvnPPgoGC2w23X0IVhhnMF2bc2OHZU/MrtQyLagaYnps02pkM
r6xXcnCZhEDfEoPtv3fLRSnA8lwBMIK4CruplZ3JrCrbwnnzUcVeDJcedmA44MgM0DQS5bR+o+Mh
B08JYKMl8aW1qZ1sALeX552INsGuM7SfQEYZzvkTyvq26ztOdazZtzGTuf9vLI14jke1NZ+pE+vT
zvU6EWtlop5gGIpVhPm6HKVKAuBQ4QJjRj1zrZZoLoYs9P5eJ3lXi0JJv8KPXY8ExTzSFHkkxrjd
o4yApQeOBV+Bq6v+aLQGDf34XsBQOM2iS2K3ZG4PWSLpj2hViuVY3k44G+zXUxEXmtMa3BkULlug
3/L+onw2K3q3gxkZ0MrafxujMs5F3AVhFYfGyHXMFo+2+CcRnk7pXD1MI+lktEHFhXnlzabeYzBf
Vtx6KS6e0lJPyQr9kBb9blkqAggDTyURb+sons4Cjl7m8y+GWf2zYlIatxWfmcjBTLuNJsS4hXZQ
OPREKszZxiX903aLzEaiJZjLKDVPxBZj8w+g0a4XoFk257xHk48M58A75//oQzzQjR59NemeWc6V
YJhyHVzVrMm7V4HS2BALqJIuML9Wy8OBBb8e9kpU9t6OmHQLwA94Ey+IyTYSsavGsDdzEB2T72Fx
n98hohb6vDpf17Qv2Mj9s9PfcgmYjXIf7xLBmJ8fQ1Ud8W0MJ2dlJT58nk45VGrgBWH6ZBPadFU2
W/nFonq+SsSt9O1W+NJTOv6i0DEy/OnV9xYAGBmZDCvO7dovNPpkRfOcvLAi91noQPNO+Ab9osHX
eNwJi8rhPr/mxc8DDeIQz8xPxBXLjC8oFPsxNm+Rdt/LZ8p9riaeYAwXuoBIavbDRR03VwvoN8gD
nUtjEe1kYBPyJHoiWuAnW23qPFWwSEUDuWc37O69VpQs88boRZyfQkBgaWEplK6OiX9EKyGirEDN
C6zvSO9sMuj5cFwz+s5a/X3OQjyaF/vq8JLag7kTFqkV3NsotcqcWnu1NNOLNWuE3Em3pCncGTWQ
J33o5Avk45Sqbo7hLJbjrLb2ntCJQRuwctp5Npm8K0ux3QZLyuTsyVPEpVdYUim8YzgdgJo3NCrp
BbXlaTnUaFCtJW161lqcx8k6nWxe0ysCSv4xe91yNB9kbiyic0CMMLl+RDycWba0oOonpWMlZESq
ikcLjrrC1JEA37kwjJMK+IFf9XQRNZnsLkZZOOLITmKU6E0vn+mP7tjOq73xNZWDi/PgpzK7AM4S
lI5Y+m/8zpvzUi7dTydtU9Yr0RZaJvIvj28TPzotDhdZPBTC35i2m5EdWu4oaK8UF/sn+O0eqPz9
m/XDOC1g9+JM6oMWQHz0lmsjY85dvKZk8LSFE2IPh2Fh2lZJpiU7Q9ttnEDgcH1AasUsOURfvV+Z
w/BxH64MZ79v5ZdfyONgObTGMv1nkjYgHhvwXV3+0aqLt81+ogRAF4lSR0lU5GFU8I9B0ULMjqHv
xLDB7wO5FC86SfJA6aReCWlffC6SuYdQCxHLMoUKRenhFBr9wNqlAyebSRsM0xXgwEhHXcgvWkV+
raQbcjBvhcmzC1lTAijkrAoChEBXxPRnV6ckFfZYA8HZOR/s/aZXcv4Ai7r5dqXX7JtftaLeX6BU
qh8AY+0Fxn/UwITUlEoAMzHPJfgMCMhIZ2bQQe+q979kudGdDm43zsphz+f60PJ+cHilKBvQ7HTN
Go5L55RN+gVVPhJeeEg0w2629PzzUQfoj7maTH1wQrHtolopqnWu9adTHNSgou791hyDYr4j14I8
5dwfsYY7S7511upjd2b3oFzO+6c+xpz7xyjgJgMV5SzF1qnoF8GyXZHYtUpFjycQ+eg3jNjFIpa9
VUwJ5vPpHAeipjXJ4mZWz9ieZV/Fweq3lKoSoosEhUw2JbWmvYihtFi0VVLYsxyNmkZInLDkln36
w8ZV/5L3G6y10BKu5Bue7RLujekjV7XY2sorC20LrxuB9dqfuS2IGq4eje47AclWGEK2rS6qzEe/
uMqAbCMYLHirfzj7SaNKPQCWJ+C5fOKbwBcwG/rhPMX29KL7kaNjqcKTvM0LzX0It+QYiMMi30uk
6dN6Zrp9rwhIGU3RVXo0tp6eubTKqtvFQeyh9QHsBcL9jLZriqPuWLKh2lbbLdDcrsJXP77h5GNH
Pf8sJR2QtW8/jHZizGiFa/VHbe8p2QzBreRTWh5ta8AuYAaod8GK8/V0vzpUCm3D1k90R7h/iYai
pfNe2BvDkHQLg1UbScCFpAHNVF3RGUHOln7hcRWCGadPQq7BFqxbIOZnecscc5DtB45c5rawE3Z9
/Rv65J28tQqelkT8REewgFM49QuddKtl1cdl8JFR1XmtKcU8lNsC2Q5/MuYnInSGGGJFbt7Xu3Jl
Sog3KoQpoeZVGGF6V9hmUP2+41XvrZCKFSZ2EPc546Y2vvhAbQw1Fb2onBcFR+n+y76iC+2Z8RIS
ecv9ZCd9RQYw3FgahFHRVrb1S0nqfnTUafRcc7kNvjuyywZJsMK2Jrt6VCg1fVilGyBGOBtUYXXP
xuv6/wQ6qUT4K94LvqVUsCrGk74RiPwSLGuHs7VL7tuu211CpIonEzvl0yw8TdCP9ov2z6Nt0DjP
jLe+ty9eyakEfgFkGx1Qik0E4R5eNPJYQFKYRNCF1SkJQddXRLiDabAJhR/o6jIZa92Q+SfDM2h8
HV75VPve+nb3AsD7GeEgoJmoQz4O/iGL/EPLqa/BBXY5qXfcQBYLNyrAsPMIEIqbudiwzmeTllv6
Af+3gtfNC2QBUKVMyqOU9i3Wix5OuK3Tww4qRrd+zrORPCr/N1bSODSn7FAppN/NikyVOANqQl0o
NOzD4g0fjg9FK1GOk0+Q2XmG3iU6fWXI3wCjx2nnvQaKDMPBj5X2ztd3iAzn4XBQnCuhavO5m1TU
c4dks9lSfndiAg/4b+1cEAiNBCka0pzwvpueH/Biu2qqYNiD9NYkwdJ1L79AjbWYIu3h6KXMQgdp
uxjzCdN3LIOD2cOHI3v8jku3FEg5jGBJurK52iAx2EB62pAtj3a/pStJZBqCFDNxN5XmpAHiuDJE
E+Wuav9a1q6boEYuOxD4aXx8nv5eG/M3ZUN5bwyqEQ5nzHTTX5cqaKpX7O1HFXbGKMoJ87bEpfLN
L7JJ/+pSBEqvObOM+JC9jBG/2PwdgcDAA4aVu0oCACV/oHMSrmi59W3A0+6v8tqrzaQ2lpd+emLE
hL+4KVNeJYru7yt9rCjphQsltGG1JmeNHOvmNxEI+HVLf1aEPAjqVs2dpDy35zlCHSvtJJNu2n4+
NkwA1mpAcffRQx0P9PJEDoFXwxk+2b8DBKYv4LJy+3FJVpzOUvcX/Heg/W7lyxWGNVEmfd8vXLTj
eiQK++425peqTYHp9gtjffxd3hRyITlyf5nJbZM5oSlPj7ypgGlkVBVlsfG+S4g85M5kVxSXzYnB
L0hF5gbjxAmIIIiiJlPL/oJhoE3tTArFYkjcPd9gjvx6F/oiLgOROcTJdsqcaDW+sLfElX5sgFty
pFnpH3LJQdzZXPw/E6te4pwEDBPqdB/u2HpfaCVFOOPd9IG4uUYwCN53Px/J8bKPOWWf1GQzgUTi
SRMlEOE66XD4PhKMxg4oe+XFecMS7ENLiSdGbI6VODBfAxcCb5GjvdTffMrm4ruVgR1anHyXm+cx
fU7iVLPeGnNEIGjgmlX5Z+FBluBKCVLmNnZC66IM99s9UJP+YOUPyvCUFun9w+IxHsPQ2y/Cs7f5
kC16da5kgDokteL5laeRIBdsHrmLet9PaljHwHEwdLcIAPK/5tG/2UTZa+zSCZ0XPWvP/tiPxMU6
L040Y8h98yiGWJ6KjiQylBNf+oOirDKwcfdgXMDvWaQ/MwxbPh+93Hx/KwwvGMUemik6uMOn2Nph
cj2xXQ/jAp15E95XvUrHzpKNJDWnnF0q0ThI18eEAJpC6V9Rir98SZWkqsW1UklMA1+TJK+H/wk7
eBS27jB9RIzEFsyAagHLk0Qi+sShEpmciUC2XwFG5/evK2WarmJbozNTgUm65pe5VD9EFrimi7EO
d7T15pc+inU0agBFUvLVpizvZvH7SA2lPYEkpAWBRdX4VZiGVgSBTRFYH3H2bPp2+f5l1uz5Dcyu
bmrWIWtR3yLDuVYp3qq37MT+6bW+MZt8GIcRPGHsMRYGhBSS+fRUtwMUfW1aKk68M3IbNUfWkANy
+dpcvmjyau/VXvHfrQpNNefnl1sJX+Tyg0RntuEy7KGSFNMIY59n2OfrHf+rU4b3k+z8DHXPNZpu
aWrPF0hUx1pnFdXz2NVfWi7fjQx6gczOuOgttgImCwmGj2saVj2bkSBxDtX9489GI3gwZMskYdeu
xCbJe0dDrjyxiPYU78Hza9sEYMrl55K6LDNmtpMp05WRDOrG5+U4wpjCn9ts3Qp24c3riUTzE+Vb
XKG+qb5A0fSbYgNnQhj3Is19b5GZdOzt2RzCAqcrPQL2V4BTAa1oOAd/9H2xNmBHXLhTPWIhHm6S
wAMYgLR99mja4ppfPRXsuWPNPcDUmf9177KuZibjMsCQZ7OhWV3i9fkpQ/EhANPbdLzxwFzJrxrq
HYDm0t23w2Fx4RayAkaUW3IWwXAGQBdnpoy6bpWMHE0Kr5qJ6pdgRkLbRfVdAmmf9DgGabaU9ClE
0h8+Y5ravT4PUEWmiqA+HsLGiVciRXoPQSIBfNgwJ5nXjyIO68yfUOgFt6czr2vcy+Bxtj7vApRJ
ALUSoaasJvIzdQCCv0dzQkBDevTtpgzKJNsaSPR4IILpYU/EatuCkh4qVtt7NyBuyIsww1E/8BW/
eIvyiYgDjJDuZkSNWRl7Y2cj+IYzzN5Tis+HvoolBZoeRgM+C82xQ3xBmfAGMCJzCcmXq2LO0ujv
Cto5kIXnHxhG33hdM7ZbTyjIc3GtaHgczDn91EVB6CzOY7kLN8+NSdjksuHp0xT34M2Sbxdt2g1x
ZWvIOXhPwrW80i0InTUpQR+p8DK4WOfxY+vHK2NPcrZ167vIFz5gf1h8UkhGUJ3zOmQ81CwdG0uf
5s5Q6VBH/kX1hvBOhBjo225w/AZfOOqaj4vw90hUpKZdYAgfVWdiG/m+Z92t13d8rTb6Rxy5Tr2+
OYQikCJ3+BAn7n12mJx63f3g8tcMmI14YObMaqPHam20DXvZWvA3H+D0J33ZIGY7pG7m9kt0ZQ+0
pNo+nSaX3aoT7ZcBLI5UZXluaZbRcrCo+1vylDt35E2aWepSL1u1sIMmWA4P4yK332pdXjm7HxA1
HumRFk/7tdVNiRL1SOd+ThwJ94MoyU048p40RI9CAXBYbBiIaNp20Z4uanS9pfe5wUd2nbXo5XWg
X1gUwpS1gSefetxxgtML0N5Od0Qr7XLwGrzoZbBSOklmYp+POJjHDVIH0tPEl0QR2D99XJH+oh//
THoB1qWZWQ+uxXMJ76bJpggKdvoFNzybn5tpoCrQ2K8Yty33E4HZTyE6YlMPnE8sBMH0fopvE1QR
oJCUtaQTBX9p/WtM8wpc8hpT7bR3wXZRmUY9F6LLRqp5NbXm5HhfDmz/9l9K5Xr10PjykWDMMNq5
mLyFNMulqLyBIF/aWw0JTvTntJniJwYGAMWgMMdHb1x4lY/WSbnq5YwEpyzJInsrs/kvy+m402UZ
p8xoTR+U6DOZieyHoqFFZuVPLWPFvDexZZ4AGsj0J1Lk0WJOA9EDlq5A93Ghi/cUkLt1MlQiOiM+
6/bReB4Ty2n/ViiGF/9yZHIZh8vVXbScuUYDA3iNw306KVFuR6MzCqHHOXN5P6v5K79SUS5/SWOE
kOijJKFF1MA3Uh5uQx1SKomxOjedpa+qWMHHif/a3zxqUjNQWcjmfTaCo8Fa8sc8lL1OHURiZDrF
WTKC3xuNpa8WXr2nrM39N8/qhTHw+xUnrdxDtdnya7wZURfEnZi3jyfiMz/7VXgd5IedF7IByhQj
vWT070usWSXobNLCn9sJYBPU2hRoKU6ba8p5ibq8znuuees4CvIACv+HhkpERExiOU7c/P+13PvU
/kcS+BAr3xux1DAAV/D7eVOyf/clitWwutGme2lBnhCI7wcGUF36gTlQqOBMVyFLdClDK+OQJdAi
IJJvdaD1tykluJUaFHRRL0pQ+FMvQwuLr2TOQY80dlDpXyCBFICQVFMPFo8U98HsFGTKP7W3YOwF
aJ8i5Uypm/G3B92hL3Sv9EVXFpBOkqYeTgPLDmKIlrI7ZCLFkbGJeHToqe/cN4y7TsjDrUE4zPKD
xdLRpkQuYYnldN6nd83Ro6+nc9kD9krsnnO6jH8zqZqbCweIu1c4gxAj0bIcWVpf32QEYYfXlOxE
xMh3Vu+c5uFLs+Kp6rie84giVdPblQkARKfpHKDbYp7U5ABvEeRrXDUSOXUnKLMiFboxJ90Mnk19
lwgAye1zMqmzzVYOAySuog2pH9nWpAbZsx7KniTpAMeZ39bjLxIhUV3ub15GWZ2kichkWUz2yZW8
0S54QwlLBWktyYFq3fV0GSVHiz/I/mTtB4OG1N/dYwvwuSKBZbGrpR83xIFaakqufO3VXLRiVBYH
vlgvxBueT6jjmEpOo5qPoeEjvWU0aWUqqlDEumkZbfFNKQq81Yk+VFJMXblODPvIe9van4d0C5Gu
C7VK6RCR4SpklklWgVxr3UjY0zoYA31PfkRLZ1XC6wvIEqO/MXzTQDdzAuFJWTtmSuNfqrd+kmlr
Ozv90tfwSxii0EdrYEEfs0etJE83Mow2dqflCLL228pYUmws3QBSNPGAVZWRS7NhfXvWAsLwqJzh
PXKP3CP98y+u3USnbNcN2qksMYnIRPFQ3IGuaQjo8LSoSyX872xduB7Xl539T6QOcbD4S+5lB00G
eVDmQ96u6JfQ+swQKtu8nbxbzJxS13Y/FVzmkShqM1y8n1+BqujqJeyD7S9LyJ5i+dxeqY5K+h9C
NfkQiCMghrEPM92Zg0GpTvkZmxq+nZRrKljC0CBLewsqopKOQc0X/7a3B08/aX3p0rgK+SGFF4lF
es2NrMfVm+yEZQl8cnNfS5wIy1SzpOng/o8MluUZTIHwrQQUgYGTaufht52JTKUV+huyFW2DAcpr
bRXZvqS6WlISD1oUZBa//+ljp8k/+Q9YVBTzEW/+eLUc4ElYBt0yn1b7pstrvGywau0apfrXbDLY
ec8HkKTVvbI1LGyo46GiqwpTRl6U5CLkhecI7BljPlN/+5yf7HwSemVC7lAwLABF12nFAX/TEkc7
l+eeJzt0Z3jMf1A3bnZpz0w7okvaXexubn78IjdAkZoYnn5+UUnf+CHS9LATt7g8e7MyUTUa5mWl
Ssvi7ILKwAdndRuyN8Sddu9J3opN4LjaNWYgoxfH3v+yw0Pcwj5NGhfY3kZp0bkH5N7gmb0ZwmaI
28miVGmqsHEjPdggxvJYEEkY+6jo3MpPaytGqBOACHrhIu8DwbQ7h57kNfOaiWwRhXl4cBGtLKTU
GX0nPSi6znk/kO8hnNm8xyr+8dcV3l9m6tPtL0RWExsvK0ZnNDZPmRpVb5IsFJlpqqcBRHXy8YyD
dmU1XzNVmobYItHu1OVPZuvZ/YK8fMKR/c/zh4P+HAWt3skawYYbRSWhaGxa5/U/jmykSaMG1jIw
x9E19zyRb4Cmk5GkGyU9jbvwaP0+pV3Hb6JWPGwMo4m8IhIMf2On2Y7uaJzcj0uIntmGAhdLxrfK
p4vqvbk+JZfx56VH1YvFKuTA3tInvgfE0J7h8mpGj5shX42sMLmF00zt6mzWjNq7ToxPS3w26Zu8
JOPvW1zUg3SUyS/a0ziZrsVgp/zksf700/nhk8Z1rJgLOHPN3ukZe2mn+1Ocr4EveE2Dj2rt1rKz
sw8FIuKfulG/FzU8LDdrKnnC4apf21cOeehi/u6yw5BKcJ/DzBSJJLkTlCsxntzTYiK3dIeb8FNu
z29vOLe8p1cmxlzz9+Fvc7oOxI6Xc7otVVwV0cKMxyKpwacYsVm8ENl6FW0uZXsrrIBzWTwDYl6e
IzREEuGFU2MbbOAyCep1FDWHWnJry/axcwK9fAekSRTHwwvfQOeaSAqotadm08sFebDa9be7bOCU
WxFvPOfQCEmguGAFP9qWKdtkpSEwphUdNLBOVjHubxxpH8zrWAAQxkX0Z+wAjozaD+VrFVWpMuNZ
6UQjd7kvWQDO2l50CYyI6Z1Nn8CPj8yfIi0xyA8+qSQqWQG5MGEIF8Qd+DM7rram2kGEutQYygJ9
gNFm/EyK+zxLPq6n2ZmVQdguwGnmcuqL/jkVbmueGeYbyAWo23wqQlCoHSV6Kfh3unTCdtV58V2Y
jW8M1dW9SHfkSSkKUluBh63oSqcSq8fRw5jqDEmN6hRtE0T+Y4cKnIxmIm+QlySiONCyfTuzhglt
hiKs5PersdPpwTpnh+C6M+RSLe7D7hY5d1ve+P45aRz3nTQ6k+9Fn7ISbh99VxIzmzIARyO0cd6O
vVI2iMSZJ6b6bJ/KMVL4NEx6iVsRQBHqnc+baTd69jqmc662VyRiMASstUEkqREjzVB3X5+w4nDU
fGt658MYn2lLo/LQbgH7l8L/KSwaHFWxhky1zPmBB7X+mtyJskUES7lELVF8cm5QQk5eX4DOy86T
tPZx508WzvRPL5FPGDKPSz3ZWvGN5DlkbS/XgVTJPxaFhceKXjyXV21JVc2aBmO18qo0J3HP3Bw3
6M+DZumyo260/uLVlcyzHk7H/tswX8/NAr0AYvKSaOBO63QExS0yR6rjw5oqo3WW632bv1xrpPw+
g9d80pGASDRoy5gzYwVcKuc4kREHvDtWv78oagiU8zwO1QDVKkc9QoDnldlyq26iZx2DUtZvgtlK
YOoHZUqtgBkT26P5zLCWUFf9oxEtakjnQX4vXp+Ts+pD9u92gwfc6ZJMeZ61WuOdZga+zqHTTh4p
fWb4FFBYcRik6lW+H9mSA/Lp58IT2CSFlRXMfk51AaNDfAFD2m3VmElRfl8rQ8A+VOYoOj6rBRao
6jjo197JNPNCZblNJkEiu3pTp/Q0upkY2pdbYAmzPhs1lXqrxwW1G//MhVey6pOjMbppoixkCvaz
NkLA9PjRIdgHW9LtHiixsvrm4wCyxxA9KNX1GnEXvkfsF/hXHbGa/3vFsZ/WIh1HxCEiaS1dIUJK
wqh2UqfydFrCV9rhkuSE/G3hLA1sT0TPrSxQ8qOJ2w6q3c59RNAWbR9MHyo1BjVGjpKZrz2yk5yO
GG1B/c1JbrYhbjmeQKbgUGugbYM2KxLo2wpipX97UlswqZmN++UqXJfvc1uxfNl/Jcl5eosY77MA
NRZ8Q/mND8fYpmzjnEWK7N3EQJqTMHxWHClrfhvGkjBGp01mYZT/c6gcdaF8JlZ7GOL5TQGT9t1e
vO/S3HH2HhlpxXb155z+cpcMxfkskUBVy1kMBdrDUR6bVGjne0ZPPLVjsZZTd088HZde9p0tsE0A
6Xcxd5cKJYc8TXlqmSpZH9dAZnT1WuhYI6H2P3zLBaYDTghMSssDf7PjCt5miASX/MdExRY1BtwE
P2n7RKCBGI9CQuadeBj2xxqW0qEGgX6z798qSWQnT6h4EqDXTv9y5IIMTm1tO5Zq8J4RnOT7rlh8
LpmT/fjZlCmOP3S7YcCqBMNrOunElRo7iJzzhG/kAQoTev/lh0C5kGq9dKYjjtTJkN2JrfX2Ohz+
1SCd5WEpo0sgi2pGXcgUOucwAvrYDGQJljjsGiLSEJzZe79mdLy48yp3gAU713vDBk+FANiIVb85
0d0g8BMmGbauYuACSsCSmzS6/TLMEyGN5JMTXRMWr6VsjOuwnZVqF5Rjsz1kLVWllpFEPywyzRc8
hae7qYaCZ11RGShTSnwp9ZpAMoUoht/YLHkknnG3PNLnw8x5HbjwVDita9BhUSQQ+Ry0Y+QRFcLQ
JkTf2TILzXnXDpz5J/vq1/U8z4i5ZmP3oDijGJlqo+GOcNIiSO4W5gww++4TqGpSZQ3kVND2ZFIY
glMA737Oh6C5dRCIQ/7qblxVgVt5S9sK5rlmIgJ1PsnpEPcD+7PFeWkmBKO1ra0ly6tUekCUuFi3
ypJ+m41oj9YVpZ+DWlDJhQHCGBRxcnOMz4B8zpns+GfbtKzIvrHM6zQpF6BXdJPi13cWpWdmWC6n
hrJRazxSG6XRWJyE+W2IB+iCa/U8CdVPb13ZJ1SPq7wWWVOOZyZeyGaLVGENyWRy5YtgSJASnleN
PNtaOqUOMOZar6cv7ybIaqAmIWXzDPnpE6evhqXpsU/1CfHrX5hZL0xMenVELpn7y+531EZb+JFC
/THfy6khTvIrsN64OJWstr/CP8hgUiMAYCLAH1o54CVZMw9z6bddy96Q86Ty6mDYtZYqXL0aV4wV
phU6aE162DdYE/tu+PJMPyMRgyW+5AZz3G7r5oWoDtD6xU5ZPc7V1PaSTfg719HJtn1tgUmWQRiH
tBq1rdzDhYTs4z4uHTBGaKuwtKkxFINSs1gUxLcuqdxJQQaRccz1OlRj+jmlxZFDMNDI5oL3gW5G
eYtgMi9lI6BZKH4A81W+R9B5FGYPZSgppkM35bQ4XLJEQqOwUVGJK8RB8RUFTXMmkazDk1/YQ9Rj
5hlbDvNp
`pragma protect end_protected

